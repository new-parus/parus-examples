netcdf in {
dimensions:
	time = 132300 ;
variables:
	short time ;
		time:units = "sec" ;
	short amplitude(time) ;

// global attributes:
		:type = "uniform timescale process" ;
		:title = "1000Hz sine + White noise.wav" ;
		:t0 = 0.f ;
		:dt = 2.267574e-05f ;
data:

 time = _ ;

 amplitude = 14, 3560, 9942, 13318, 16720, 20263, 22867, 24907, 27126, 30818, 
    31749, 31074, 30233, 28827, 27869, 24764, 23035, 20892, 17196, 12402, 
    8741, 5325, -295, -5194, -8058, -13583, -17666, -20167, -23609, -26085, 
    -28522, -31121, -32098, -31684, -29179, -29775, -28855, -26747, -24670, 
    -20525, -15219, -13161, -9129, -6499, -1011, 5147, 7707, 13162, 16748, 
    20224, 22817, 24826, 28495, 29671, 30916, 32054, 29099, 30081, 28338, 
    26194, 24086, 19072, 15720, 12022, 9262, 5633, 1165, -3048, -8369, 
    -12054, -15445, -21099, -23980, -25253, -28109, -27828, -29597, -30825, 
    -30246, -29282, -28480, -26178, -24163, -22345, -16219, -13549, -8705, 
    -5602, -220, 1988, 8268, 12172, 16192, 18787, 22988, 27063, 28372, 29233, 
    29201, 31367, 30306, 29250, 28401, 25511, 25238, 20827, 17466, 15034, 
    9688, 5388, 2039, -3564, -9008, -12623, -14750, -19480, -21684, -25242, 
    -27183, -29821, -29031, -28911, -32004, -29222, -30234, -26692, -25753, 
    -20669, -19154, -14634, -9470, -4551, -1410, 3219, 7096, 11412, 14217, 
    19595, 22931, 25717, 28343, 28711, 29955, 31044, 30046, 30414, 29579, 
    26675, 23552, 21576, 18911, 14045, 10825, 5516, 2705, -3303, -5958, 
    -9746, -13535, -19186, -23142, -26033, -25718, -29022, -31275, -31350, 
    -29923, -30620, -30461, -26916, -23141, -20946, -18312, -13042, -9460, 
    -6080, -2679, 2137, 7842, 10688, 15173, 19564, 22836, 25396, 28356, 
    29188, 29128, 31581, 29169, 30159, 27180, 27366, 22689, 20775, 18814, 
    15408, 9850, 6469, 2163, -2468, -7583, -11129, -15270, -18399, -21423, 
    -24942, -26063, -28069, -29691, -31326, -30863, -31024, -30148, -27471, 
    -25065, -21141, -17494, -14334, -10356, -5830, -1466, 2896, 5877, 10203, 
    14343, 18544, 23105, 25868, 26578, 30182, 28943, 30683, 31593, 30170, 
    28369, 27916, 23999, 21379, 17320, 13659, 9409, 6240, 1517, -2765, -7583, 
    -12015, -15270, -18634, -21178, -25433, -26550, -29434, -30698, -29751, 
    -30638, -28683, -27816, -27139, -24620, -23215, -18540, -15072, -11570, 
    -7216, -1998, 1994, 6361, 11722, 14296, 18798, 21515, 25651, 26494, 
    29591, 29718, 31235, 30499, 31836, 28903, 28122, 24896, 21050, 18467, 
    16022, 10607, 7585, 3073, -1861, -7025, -8841, -12757, -16786, -21323, 
    -23068, -25311, -28908, -30140, -30464, -30945, -29145, -28419, -27266, 
    -25422, -21751, -20019, -14532, -10651, -7626, -3794, 366, 4880, 9544, 
    13545, 16200, 21562, 23193, 26064, 27055, 28969, 31292, 31024, 30373, 
    30229, 27419, 24526, 22323, 18604, 15865, 11413, 7315, 3134, -1927, 
    -5758, -9480, -13712, -17048, -21522, -23032, -26518, -27058, -28989, 
    -30059, -31520, -30968, -29434, -26959, -25485, -24160, -20328, -17166, 
    -11970, -6479, -4266, 1397, 6467, 10126, 12209, 18180, 20875, 23385, 
    27756, 28768, 29737, 31084, 29671, 31789, 28867, 28504, 26997, 22837, 
    19569, 16242, 12313, 8374, 3729, 754, -4047, -10945, -12808, -18121, 
    -21375, -23193, -25724, -29529, -30123, -29614, -30548, -31365, -28796, 
    -28478, -24934, -22785, -19300, -16145, -12535, -7943, -3749, 689, 5276, 
    10433, 13310, 16455, 20511, 22196, 24772, 28477, 29018, 29807, 30191, 
    30483, 30569, 28772, 24688, 22573, 18104, 17918, 13719, 8151, 4428, 445, 
    -4682, -8651, -12780, -16381, -20114, -22873, -26801, -28366, -29735, 
    -29365, -29436, -32312, -29435, -27560, -24467, -21923, -20330, -16223, 
    -13588, -8597, -3222, 569, 4569, 8802, 11901, 17601, 20185, 23896, 25656, 
    26884, 29001, 29718, 29800, 31070, 29022, 28780, 25790, 22849, 21942, 
    16669, 12873, 9591, 5345, 1090, -3910, -8144, -13165, -15420, -20638, 
    -24367, -26312, -28557, -30638, -29744, -30318, -29662, -28752, -27548, 
    -26252, -22555, -21305, -18247, -13242, -8885, -4500, 826, 3208, 7585, 
    12899, 16779, 18831, 22777, 25967, 29159, 30344, 29996, 30189, 30836, 
    30705, 26608, 26915, 24804, 20735, 17568, 13900, 10482, 5749, 14, -2289, 
    -8118, -11202, -16613, -18524, -23266, -25581, -28389, -28798, -30927, 
    -30150, -29956, -29976, -28762, -27520, -23129, -19621, -17738, -13196, 
    -9530, -5035, 604, 2988, 7506, 11460, 15643, 20499, 23276, 24119, 26441, 
    30808, 29880, 30558, 30873, 30668, 29236, 28002, 23531, 20634, 17688, 
    14029, 9708, 6080, 2182, -2433, -7281, -10995, -14059, -18696, -22587, 
    -25760, -27514, -29562, -30941, -30825, -30798, -28710, -28048, -26347, 
    -22754, -19651, -17577, -14302, -8406, -4892, -2129, 3893, 7386, 9833, 
    14548, 20347, 22681, 25116, 27363, 29190, 29331, 31823, 29239, 30583, 
    28450, 27280, 25033, 22008, 17467, 14598, 11097, 5598, 2924, -3342, 
    -7787, -11757, -15281, -19570, -22140, -25324, -27724, -29351, -30084, 
    -32303, -30844, -31081, -28546, -25928, -24905, -21248, -17838, -14527, 
    -11532, -6435, -1876, 2677, 7240, 12334, 13941, 17357, 22499, 24351, 
    26924, 28826, 29239, 30612, 31089, 29114, 28726, 25494, 25773, 21952, 
    18001, 14090, 11227, 7320, 1249, -3004, -7520, -10189, -13811, -19052, 
    -21965, -25826, -26437, -28944, -29994, -30109, -30592, -31561, -28558, 
    -25760, -26027, -22334, -19721, -15211, -11483, -6711, -2670, 2679, 7026, 
    10101, 15300, 18767, 21857, 23956, 27323, 28914, 31133, 30278, 29229, 
    31205, 28004, 27654, 24772, 22139, 17842, 14279, 12020, 6922, 1000, 
    -1473, -4500, -9120, -12811, -19069, -22380, -24530, -26217, -27814, 
    -31269, -30802, -31687, -30134, -28391, -28868, -24109, -21984, -20270, 
    -14181, -11007, -7833, -2570, 1747, 6838, 10106, 15736, 18785, 20126, 
    23401, 27235, 28955, 30580, 30045, 30769, 29715, 29043, 28803, 25509, 
    22570, 19011, 14239, 11452, 8356, 1845, -2495, -5691, -9205, -14179, 
    -16997, -20631, -25031, -27285, -28676, -29618, -31004, -30905, -30519, 
    -27990, -28100, -25757, -22065, -19190, -16846, -12135, -6440, -3901, 
    1061, 4678, 11150, 13784, 17598, 21005, 23216, 28073, 26895, 29523, 
    31149, 30850, 31225, 28949, 28407, 25669, 22635, 18953, 15509, 11293, 
    5955, 3338, -2012, -5164, -8816, -13979, -18943, -19680, -23074, -26361, 
    -28901, -30015, -29952, -30148, -29170, -30847, -27942, -24627, -23500, 
    -20384, -14750, -11619, -8949, -2622, -142, 5400, 8582, 12750, 16606, 
    20576, 24345, 26176, 28429, 30647, 30846, 30572, 30865, 29567, 28746, 
    25857, 23616, 19466, 17080, 12684, 6857, 2699, -482, -5532, -10311, 
    -13912, -16596, -19982, -22047, -25679, -27970, -28257, -30900, -31392, 
    -30009, -29004, -27904, -25029, -23034, -20309, -17080, -12380, -8378, 
    -3429, -595, 3892, 10145, 11937, 17028, 20126, 23106, 25876, 28612, 
    29328, 31481, 31124, 31325, 29898, 26959, 26124, 22917, 21564, 15710, 
    11235, 8245, 3754, -123, -2931, -9244, -13822, -17025, -19549, -23657, 
    -25041, -27645, -29978, -29357, -32124, -30509, -29329, -27798, -27159, 
    -22156, -20184, -16561, -12153, -8332, -4247, 638, 2777, 8615, 12886, 
    18035, 21004, 23183, 24880, 27970, 30332, 29624, 31301, 30310, 29707, 
    28006, 25953, 23390, 21782, 17406, 13004, 7136, 5956, -717, -3587, -7427, 
    -12473, -16613, -18348, -23001, -25964, -26794, -31253, -31005, -30958, 
    -29634, -29746, -29591, -26415, -22889, -21181, -16135, -12024, -10539, 
    -6494, -616, 4347, 8344, 11596, 16356, 20936, 23791, 26371, 26745, 29078, 
    31936, 30381, 30814, 28748, 27978, 27590, 24656, 21607, 17362, 13087, 
    9704, 4587, 241, -3934, -8954, -12694, -16286, -19337, -23554, -26650, 
    -28355, -30784, -31207, -29888, -30433, -29011, -28123, -24855, -22127, 
    -20080, -17184, -11857, -10637, -6358, 513, 3949, 6642, 11559, 15071, 
    19560, 22917, 25352, 28378, 29328, 29747, 30503, 29527, 31325, 28015, 
    27267, 23669, 20871, 18231, 14515, 10922, 6013, 1039, -2328, -8964, 
    -11478, -15845, -20236, -23485, -25170, -27348, -28983, -30002, -31157, 
    -31467, -29180, -29473, -27607, -23945, -20986, -18034, -14004, -10008, 
    -6042, -1392, 2347, 7694, 13048, 16426, 19591, 23945, 25620, 26942, 
    29282, 29487, 30793, 30052, 29010, 28323, 27292, 24514, 20380, 16849, 
    13630, 10703, 5531, 449, -3464, -8126, -11909, -16578, -19408, -21904, 
    -25112, -28562, -29478, -30077, -30752, -30367, -28853, -29027, -26144, 
    -23254, -22268, -18713, -13849, -10597, -6020, -1098, 3956, 6845, 11611, 
    16062, 19753, 22380, 25127, 27144, 28580, 30178, 30723, 30318, 29500, 
    27496, 28248, 24381, 22109, 17671, 16071, 12004, 5549, 1934, -1899, 
    -6252, -12289, -14598, -18342, -21690, -24194, -27737, -27480, -31357, 
    -31814, -31785, -30507, -28886, -26761, -24908, -21435, -18459, -14199, 
    -10223, -7515, -1085, 1018, 7436, 9675, 14275, 18832, 21231, 26153, 
    28853, 28998, 29575, 31032, 30943, 28630, 29184, 26490, 24342, 21143, 
    18519, 15363, 10724, 8000, 3761, -2994, -6113, -11284, -16094, -18766, 
    -21162, -24771, -26337, -27825, -29941, -29369, -30555, -30827, -28575, 
    -27049, -26384, -20550, -17581, -14893, -10032, -7689, -3231, 1984, 6069, 
    10200, 15117, 19296, 20618, 23587, 26690, 26858, 29840, 30284, 29464, 
    30504, 28775, 26763, 26016, 22393, 19150, 15694, 10332, 6292, 2235, 
    -1573, -4131, -9676, -14170, -18342, -19839, -25367, -27321, -28493, 
    -31161, -30552, -30313, -29009, -29807, -27843, -24272, -22383, -19811, 
    -14531, -10771, -6971, -2883, 1085, 4581, 9820, 13345, 16797, 20556, 
    23837, 26629, 28292, 29102, 30646, 31592, 30191, 28801, 29015, 23881, 
    23784, 17702, 15354, 10789, 7845, 2226, -1901, -4870, -10631, -14757, 
    -18458, -20784, -24368, -27555, -27932, -30061, -30580, -31526, -29717, 
    -30103, -28175, -25118, -23160, -19605, -16601, -11519, -7169, -2893, 
    1869, 4047, 9006, 13947, 16403, 21246, 24383, 25162, 29034, 30048, 29593, 
    30878, 30928, 30496, 26417, 24291, 22290, 20225, 16897, 10551, 9511, 
    3877, -1201, -4936, -10783, -14445, -17019, -21782, -24198, -26222, 
    -29013, -29308, -30070, -31659, -29049, -28542, -28470, -25681, -21364, 
    -19060, -16657, -12742, -8104, -4784, 1348, 4125, 8128, 14238, 17243, 
    20972, 23916, 26894, 28705, 28573, 30539, 30663, 29744, 28779, 28150, 
    25144, 23353, 18672, 15426, 12004, 9438, 4380, 1061, -4560, -7297, 
    -13751, -17203, -20621, -22372, -25979, -29816, -28412, -29478, -31654, 
    -32063, -30061, -28413, -26696, -23121, -20075, -17162, -12098, -8631, 
    -4299, -1038, 3864, 8876, 14607, 18057, 19340, 24266, 26610, 27123, 
    29162, 29687, 30541, 29805, 30052, 27302, 26177, 22631, 20841, 15561, 
    14726, 8719, 5104, 1197, -4116, -7420, -11467, -17328, -20835, -24425, 
    -24848, -28560, -30955, -31830, -31247, -29992, -28852, -29164, -25764, 
    -22807, -20868, -17599, -14335, -10086, -4946, -822, 3974, 7401, 11332, 
    16417, 20026, 24009, 23961, 27909, 28691, 29574, 31775, 30889, 30677, 
    28505, 27073, 24153, 21546, 16815, 14104, 8679, 4624, 482, -3078, -7359, 
    -11134, -14780, -18512, -24276, -26110, -27034, -28952, -30369, -30577, 
    -30417, -29183, -28326, -26252, -23029, -20759, -16681, -14426, -10504, 
    -4782, -1894, 2750, 6428, 12177, 15237, 21366, 21352, 23995, 26041, 
    28902, 30777, 30586, 31049, 29902, 28454, 27077, 23049, 21881, 17917, 
    15031, 9605, 6808, 2181, -1402, -8629, -12480, -14309, -18737, -22001, 
    -25343, -26757, -28541, -31683, -32312, -31549, -29787, -28958, -27266, 
    -23959, -21554, -17026, -14285, -10976, -5092, -1247, 3217, 7429, 12683, 
    15201, 18142, 22353, 25594, 27982, 28927, 30888, 32305, 31664, 28737, 
    28995, 27963, 24679, 20803, 18717, 13988, 10959, 5103, 2282, -1394, 
    -7636, -13024, -13510, -19485, -22675, -25185, -27573, -27544, -30732, 
    -30632, -30061, -30071, -27731, -27701, -22911, -21638, -16697, -14645, 
    -8894, -5952, -3361, 2258, 6205, 10810, 14481, 18429, 21428, 24939, 
    28544, 29018, 30789, 30074, 30344, 30275, 28317, 26843, 24424, 21756, 
    17706, 13701, 9129, 7158, 1109, -2283, -7148, -10201, -14033, -19323, 
    -22079, -25274, -28662, -28518, -31047, -29865, -31333, -31048, -28810, 
    -26896, -24099, -20270, -18715, -15248, -11118, -6131, -2021, 658, 7419, 
    11380, 15719, 19113, 20258, 24334, 26157, 29904, 30718, 31655, 30857, 
    31736, 29175, 27888, 23934, 21339, 18776, 13985, 10276, 6461, 2792, 
    -3068, -4923, -9780, -13861, -17807, -22048, -24376, -28106, -28952, 
    -30455, -30554, -31031, -30863, -29090, -27714, -25563, -22368, -17757, 
    -15485, -10692, -7405, -3455, 2937, 5598, 10617, 13128, 17888, 20946, 
    24999, 27926, 27752, 31678, 31312, 31163, 31606, 29123, 26384, 25471, 
    22730, 18045, 15711, 11565, 7936, 2588, -1952, -6141, -11467, -15617, 
    -18336, -21045, -24917, -26809, -27526, -30585, -31586, -32166, -30559, 
    -29167, -26502, -26015, -22396, -18404, -15544, -12650, -7668, -3283, 
    1140, 6473, 9335, 14045, 16970, 22567, 23250, 26984, 28095, 28600, 29808, 
    30436, 30433, 29705, 27256, 23864, 21446, 19386, 16505, 11096, 6388, 
    2869, -155, -5229, -10510, -13971, -17858, -20772, -24405, -27099, 
    -26926, -29399, -28875, -31522, -30591, -29257, -26875, -26346, -23732, 
    -20871, -16080, -11712, -8158, -2849, 924, 5061, 10095, 13392, 16612, 
    21126, 23703, 27960, 30119, 30202, 30608, 31664, 31141, 29605, 28152, 
    25165, 23626, 20254, 15685, 13432, 9182, 3359, -2325, -5103, -9552, 
    -14640, -16530, -21581, -22887, -25966, -27476, -29726, -32079, -29918, 
    -29790, -29483, -26751, -25785, -23517, -20793, -16449, -11261, -7533, 
    -4657, 477, 6032, 10000, 12340, 17857, 20676, 22823, 27257, 27945, 29808, 
    29736, 30208, 31101, 30914, 27279, 25947, 23030, 18478, 16760, 13292, 
    9829, 4485, 63, -3847, -9542, -13051, -16166, -20360, -23115, -24337, 
    -28980, -30808, -31211, -31276, -30628, -30651, -29218, -26311, -23279, 
    -21193, -17294, -11751, -8125, -4380, 94, 4707, 8542, 13144, 15076, 
    20655, 23096, 25877, 28941, 30065, 30435, 30995, 31182, 29369, 28845, 
    25178, 24202, 20451, 15855, 13709, 9685, 4424, 106, -5209, -8945, -12366, 
    -15312, -20516, -23423, -25179, -27271, -28115, -29868, -30519, -31356, 
    -29676, -28598, -25905, -22533, -19633, -17814, -13173, -9054, -4778, 
    -448, 4518, 7194, 11587, 15248, 20205, 23377, 24281, 26816, 30278, 30123, 
    32192, 30739, 29379, 28536, 25856, 22367, 21658, 18784, 12632, 10024, 
    3433, 836, -2367, -9252, -10893, -16457, -19155, -22759, -24318, -28696, 
    -29158, -30333, -31115, -30320, -31048, -28122, -27820, -24543, -19204, 
    -17367, -14116, -9559, -4787, -1063, 4794, 8509, 12218, 15908, 20068, 
    24327, 24524, 28671, 28793, 30186, 29786, 31808, 31328, 29631, 26481, 
    23688, 21697, 18780, 14304, 9414, 5733, 1173, -2994, -9311, -11371, 
    -14295, -19998, -22300, -25047, -26229, -29023, -30812, -31990, -30733, 
    -31580, -28903, -27027, -25061, -22494, -17592, -13293, -8917, -6630, 
    -1047, 3656, 8911, 12050, 15692, 18176, 23614, 24133, 27134, 28771, 
    29738, 31377, 31174, 30087, 27545, 27545, 24195, 21310, 18437, 14867, 
    10384, 5381, 2832, -4292, -7930, -11281, -15574, -19589, -23688, -26046, 
    -26618, -29103, -30961, -30499, -30393, -28939, -27205, -28234, -24901, 
    -20218, -19181, -13456, -8800, -5887, -1185, 2320, 6550, 10952, 16586, 
    20286, 22318, 25060, 26433, 29894, 28612, 32574, 31363, 30515, 28834, 
    27872, 25168, 22831, 18118, 14724, 9995, 6635, 1152, -1530, -6953, -9227, 
    -14719, -19237, -21894, -25294, -27457, -29136, -30106, -31706, -31335, 
    -30696, -29664, -25529, -25465, -23082, -19113, -14160, -10285, -5400, 
    -2458, 1184, 6710, 11839, 14045, 19044, 21110, 24646, 27158, 29287, 
    29864, 31766, 29812, 29423, 28936, 26247, 24717, 22356, 19440, 14834, 
    11363, 6898, 2665, -967, -7059, -9829, -14655, -18014, -21915, -24500, 
    -27822, -29437, -29836, -28983, -30516, -28856, -28187, -27199, -24805, 
    -22235, -18132, -14728, -11342, -8261, -3309, 1232, 7323, 10682, 13832, 
    19214, 21790, 23577, 28055, 29729, 30135, 30805, 30823, 30124, 28268, 
    26483, 24402, 22829, 18538, 16439, 11320, 8332, 3317, -2166, -5985, 
    -9683, -13121, -17909, -20965, -24286, -25733, -27791, -29309, -31768, 
    -30424, -29301, -27819, -26629, -25793, -22116, -18945, -15739, -10650, 
    -7424, -3189, 1065, 7292, 11268, 15329, 17694, 20562, 23677, 25352, 
    27956, 30896, 31316, 29862, 31201, 30370, 28389, 25681, 23299, 18304, 
    16388, 10951, 7617, 3107, -2167, -5005, -9060, -12801, -17794, -20297, 
    -23746, -25885, -28463, -30774, -31572, -30754, -31184, -28444, -28101, 
    -25355, -23240, -19125, -15207, -11898, -6877, -2742, 1244, 6580, 10342, 
    11853, 18062, 22202, 25172, 27186, 29665, 29783, 30523, 30393, 30347, 
    29828, 27962, 23907, 21305, 20665, 15604, 12022, 6583, 2772, -153, -6186, 
    -8563, -14452, -15665, -21966, -24377, -26429, -28430, -30014, -30726, 
    -30268, -30138, -28356, -28362, -25580, -22976, -20009, -16876, -13008, 
    -8331, -4454, 351, 5783, 9463, 13831, 17407, 20688, 23487, 24759, 29069, 
    28935, 30190, 31086, 31609, 30812, 26818, 25157, 22550, 20371, 17332, 
    12929, 6829, 5800, 1297, -4297, -8187, -14383, -17178, -20264, -22843, 
    -25716, -27359, -28653, -30733, -31095, -29727, -28312, -27868, -25863, 
    -22645, -20549, -17624, -13361, -10047, -4063, 283, 3311, 8884, 11184, 
    15997, 20185, 23059, 27154, 28779, 29232, 31476, 31951, 30777, 30150, 
    29480, 25678, 22872, 21564, 15189, 13863, 7732, 4418, 286, -4463, -8841, 
    -14113, -15538, -18880, -23643, -25608, -28400, -29480, -30876, -29905, 
    -30088, -30233, -26915, -25257, -23424, -21376, -16760, -13712, -10040, 
    -5808, -593, 5654, 8724, 13041, 16758, 20527, 23435, 25708, 26131, 29888, 
    31244, 30300, 31353, 29064, 28500, 25791, 22787, 20867, 17669, 13747, 
    9802, 5906, -794, -3379, -8475, -12994, -14622, -19407, -23136, -25583, 
    -27776, -30283, -31177, -30956, -30647, -30585, -28138, -27258, -22758, 
    -21555, -17995, -14655, -9777, -5084, 775, 4130, 7709, 13042, 14518, 
    17794, 22384, 25901, 28237, 27561, 29548, 29798, 30915, 30811, 29932, 
    27793, 24024, 21053, 17708, 12484, 9771, 4008, 64, -4067, -6540, -13004, 
    -15669, -20060, -23178, -25078, -28187, -29863, -29999, -30472, -31368, 
    -29769, -29745, -25649, -24846, -19730, -18323, -13644, -10564, -4658, 
    -1515, 1706, 9194, 10573, 15915, 17982, 22419, 26305, 27610, 28571, 
    30800, 29619, 30304, 30084, 29725, 27519, 23673, 22870, 18166, 14685, 
    8823, 4269, 1287, -3883, -6908, -12347, -14159, -18747, -21944, -24397, 
    -27449, -30613, -29941, -30643, -30621, -30336, -28957, -27721, -24408, 
    -21578, -18755, -14135, -10445, -6084, -1496, 2363, 7277, 10104, 15996, 
    17169, 21269, 24244, 25951, 29532, 28906, 30586, 30651, 29103, 28481, 
    26823, 25292, 22195, 17921, 13458, 10588, 6129, 3751, -2466, -5801, 
    -11214, -14678, -18594, -22716, -26079, -27032, -28011, -30585, -30828, 
    -31301, -29882, -29839, -27502, -25931, -22480, -18037, -13852, -11291, 
    -7437, -1764, 1951, 7395, 10326, 15198, 20038, 21308, 24863, 28264, 
    30566, 30789, 31124, 29944, 29927, 28269, 28051, 24299, 20314, 18881, 
    14548, 10909, 5934, 766, -442, -5424, -10244, -13235, -18377, -21781, 
    -25116, -27500, -29726, -31453, -30860, -31883, -31894, -28276, -28013, 
    -24511, -21785, -20492, -14924, -10820, -5435, -3327, 1871, 5635, 10316, 
    14441, 19077, 21013, 24431, 26777, 28560, 30828, 30487, 30745, 30165, 
    28924, 28053, 25893, 24002, 18873, 15267, 10409, 7187, 4524, -2507, 
    -4788, -9480, -15038, -17081, -20143, -22964, -28292, -28586, -29637, 
    -30980, -29625, -29887, -30483, -29049, -24133, -23949, -19033, -15053, 
    -12613, -7738, -1763, 880, 4480, 11299, 13612, 17963, 21473, 24272, 
    25191, 27455, 29525, 29572, 29949, 29835, 27763, 27247, 25586, 21788, 
    19645, 15996, 13009, 7046, 4011, -1566, -6554, -9745, -13889, -18912, 
    -20161, -22601, -26100, -28481, -29545, -30292, -32031, -28945, -29245, 
    -27110, -25309, -22662, -19524, -14727, -13285, -6895, -3300, 1981, 4741, 
    10170, 13482, 17564, 20757, 22829, 25514, 28598, 30295, 29282, 31370, 
    31945, 30467, 28473, 24213, 23875, 20714, 15634, 12263, 7557, 4087, -272, 
    -4927, -10637, -12884, -17435, -20736, -24093, -25333, -28027, -29845, 
    -29621, -29937, -28889, -29227, -27464, -26842, -24338, -20893, -15209, 
    -11506, -9160, -2517, -623, 4790, 10023, 13220, 16965, 19453, 22768, 
    26077, 28393, 29955, 30369, 30628, 30887, 30396, 27601, 26907, 23825, 
    18617, 16302, 14164, 6996, 3810, -20, -5148, -8972, -12550, -17118, 
    -20765, -22557, -25783, -28009, -28354, -30932, -31312, -31241, -30017, 
    -27558, -26100, -23509, -21012, -16989, -13645, -9403, -3266, -78, 5121, 
    8793, 11312, 17935, 19903, 22088, 24878, 27121, 28142, 28890, 30663, 
    29546, 30154, 28913, 26070, 23912, 21186, 15880, 14726, 8189, 5380, -146, 
    -4581, -7480, -13080, -16496, -19180, -22194, -24377, -27668, -31327, 
    -29498, -31438, -31135, -29072, -28105, -25635, -23394, -21114, -16814, 
    -12686, -9254, -5135, -610, 4671, 8821, 11854, 17226, 19099, 24137, 
    26356, 29497, 28489, 30620, 31468, 30604, 29642, 28897, 24620, 23037, 
    20541, 17561, 14045, 8894, 5115, 461, -3448, -8388, -13155, -15141, 
    -21307, -21619, -25170, -27299, -28227, -29841, -30193, -31086, -29076, 
    -29138, -26652, -23916, -20983, -16818, -12301, -10470, -5900, -931, 
    4406, 8423, 12822, 15867, 20554, 21910, 26271, 29214, 29597, 29986, 
    31033, 29340, 31121, 26771, 27715, 23616, 21948, 17535, 14312, 11084, 
    5294, 1233, -4395, -7536, -11225, -15278, -20460, -23031, -26525, -27431, 
    -29195, -31088, -30399, -29978, -30196, -28464, -26885, -23819, -20450, 
    -18636, -14537, -8778, -6447, -1437, 2678, 6580, 11381, 16343, 18452, 
    22652, 25263, 26004, 29100, 29342, 31604, 29260, 30168, 28695, 26159, 
    24373, 21675, 17458, 13442, 10353, 4164, 3163, -2816, -6432, -11116, 
    -14198, -18866, -22411, -26254, -28529, -29126, -30303, -30822, -31988, 
    -28664, -30339, -26705, -23260, -21393, -19920, -13759, -9598, -6438, 
    -269, 1712, 7143, 10653, 13427, 18269, 21463, 24437, 26696, 29226, 30532, 
    29926, 30005, 29485, 28154, 26023, 26231, 23214, 18934, 15714, 12010, 
    6816, 1837, -2932, -7321, -10680, -14596, -19946, -21598, -23373, -27262, 
    -30566, -30169, -31319, -30712, -29475, -29355, -27954, -23007, -20481, 
    -17172, -14449, -11197, -6301, -1476, 3943, 7008, 10413, 13697, 18002, 
    22995, 24349, 28283, 30182, 31824, 30318, 32315, 28890, 28647, 27195, 
    26079, 21944, 19470, 14736, 11738, 6443, 3300, -3261, -4858, -10325, 
    -16027, -19121, -21405, -24211, -26879, -28193, -29695, -30699, -30706, 
    -30383, -27862, -27437, -24118, -21866, -18802, -14483, -11665, -7757, 
    -2318, 1996, 7119, 9015, 13743, 18108, 21832, 25441, 25786, 28904, 30154, 
    30046, 30789, 30374, 28923, 28705, 25596, 22315, 19587, 14769, 12654, 
    7853, 2512, -2009, -5453, -8460, -12618, -16504, -21060, -25695, -26674, 
    -28804, -28991, -28959, -30655, -29723, -28595, -28368, -24223, -23128, 
    -19769, -16102, -10536, -7068, -2418, 1239, 5507, 8673, 12883, 17300, 
    21302, 24107, 27367, 27009, 30691, 29475, 31469, 31010, 29149, 27680, 
    24040, 21543, 19749, 14638, 10827, 7744, 2132, -1001, -4368, -9063, 
    -14628, -18381, -22024, -24389, -25576, -28989, -30653, -29986, -30338, 
    -30832, -29743, -29026, -25947, -23102, -19495, -16014, -12844, -8205, 
    -3686, 1023, 5378, 8619, 13710, 17627, 20653, 23828, 26243, 28585, 30625, 
    30096, 30045, 28980, 30733, 27581, 26091, 21944, 20668, 16451, 13320, 
    7546, 3592, -383, -4104, -10309, -12173, -15903, -22559, -24072, -26179, 
    -28312, -28023, -31177, -30317, -29467, -28282, -27386, -26394, -24343, 
    -18867, -17326, -12282, -9281, -4902, -1224, 5227, 9432, 14418, 17369, 
    19267, 22494, 26510, 27742, 29701, 30098, 30402, 31060, 29838, 26485, 
    25894, 21415, 21207, 16305, 13013, 8260, 3547, 359, -4120, -9234, -11337, 
    -16694, -20574, -24351, -25702, -29343, -28925, -30999, -30142, -30844, 
    -29605, -28236, -26539, -22493, -19683, -16721, -11775, -8914, -4546, 
    1371, 4015, 9102, 12251, 17068, 18442, 22554, 25715, 28733, 28580, 29181, 
    29623, 30474, 29855, 28222, 25609, 22873, 21608, 15917, 13437, 8712, 
    5356, 898, -4644, -8825, -12484, -16725, -18891, -21452, -24876, -26538, 
    -29351, -31234, -30973, -30255, -30443, -29350, -25571, -23326, -20675, 
    -17384, -11507, -9192, -6082, 1030, 3927, 8329, 12347, 15365, 20730, 
    23203, 26131, 26720, 30627, 28994, 31674, 30887, 30062, 27742, 26241, 
    23745, 20407, 16244, 12351, 9168, 4835, 1970, -3192, -8100, -12370, 
    -15418, -19342, -23081, -25705, -26691, -28441, -29964, -30869, -31099, 
    -29484, -27629, -25425, -25307, -21827, -17132, -12966, -9403, -6205, 
    -671, 2900, 7570, 12740, 15977, 19086, 21795, 26064, 28862, 29599, 31153, 
    31448, 31064, 29331, 29054, 27726, 24440, 20592, 16484, 13958, 8596, 
    6603, 943, -3247, -6298, -12567, -15700, -19291, -21009, -25784, -27108, 
    -30360, -30623, -30305, -30335, -30695, -27638, -28047, -24000, -21358, 
    -16487, -13773, -9958, -4973, -2322, 2247, 7467, 12214, 16737, 20501, 
    22539, 26258, 28269, 29871, 30878, 31357, 30412, 29376, 27696, 26568, 
    22715, 21647, 18391, 15373, 11194, 6904, 525, -3974, -7521, -10878, 
    -14803, -18351, -22466, -24799, -27320, -27210, -30124, -30393, -29713, 
    -29638, -27320, -27281, -24762, -22959, -19450, -12704, -9051, -6716, 
    -1022, 4048, 6869, 9896, 13671, 18646, 21391, 24136, 28021, 29273, 29574, 
    30239, 30139, 29725, 27676, 26618, 25038, 20863, 18461, 13992, 11027, 
    5112, 3369, -2089, -6461, -12692, -15010, -19788, -21761, -23704, -27671, 
    -29083, -30820, -29658, -29988, -31379, -29462, -26548, -22850, -22096, 
    -19200, -13259, -11434, -7793, -2871, 2243, 6178, 10176, 14315, 18458, 
    21566, 25051, 27744, 28643, 29443, 31200, 30067, 31919, 28817, 27959, 
    24445, 21899, 19056, 16304, 11191, 6965, 2317, -1979, -7628, -11703, 
    -13492, -18755, -22912, -24419, -26441, -28509, -29607, -30996, -31455, 
    -29998, -30319, -27828, -24863, -21972, -19296, -14114, -10497, -8189, 
    -2860, 2392, 6339, 11633, 15567, 17530, 21327, 23901, 27227, 27278, 
    29558, 29552, 30754, 31573, 29120, 26994, 26479, 21502, 17677, 15148, 
    11354, 5921, 3187, -1065, -6215, -10009, -14016, -18274, -20027, -24161, 
    -27187, -29540, -30847, -31644, -31065, -29408, -30106, -28903, -23992, 
    -20823, -20343, -15601, -11625, -8041, -4092, 112, 5390, 9028, 14079, 
    18080, 20762, 23183, 25631, 27637, 31155, 31341, 31280, 29393, 28617, 
    27693, 26079, 21007, 19062, 15038, 12354, 6815, 4322, -886, -4406, 
    -11466, -13870, -16517, -20909, -23862, -25187, -28721, -30632, -31115, 
    -29776, -31617, -30372, -26948, -26315, -23018, -18834, -16959, -11371, 
    -6578, -2539, 1819, 6194, 8463, 14231, 17074, 20270, 23346, 28010, 27871, 
    30783, 30592, 30398, 31968, 28839, 27090, 24772, 21791, 19587, 16216, 
    12479, 8190, 4797, -1204, -4871, -9722, -12661, -15961, -20614, -23490, 
    -25450, -27653, -30671, -31862, -30643, -29379, -29923, -28397, -25082, 
    -23421, -20061, -16027, -12046, -9343, -5301, 259, 4239, 8980, 14247, 
    17226, 20513, 22387, 28020, 29448, 28532, 28826, 31126, 30717, 29852, 
    27507, 26007, 24129, 20348, 17633, 11099, 9427, 4383, -408, -2797, -9743, 
    -13809, -15539, -20215, -23667, -26254, -26584, -29339, -30683, -29640, 
    -30380, -30932, -28220, -24090, -23366, -20439, -15213, -13533, -8678, 
    -4654, 101, 6064, 8956, 11238, 16149, 19951, 22724, 25114, 28711, 29911, 
    30761, 29259, 30875, 30698, 28862, 26141, 23645, 20310, 15574, 13687, 
    7649, 4955, -303, -3662, -9055, -12936, -14942, -20767, -23892, -26475, 
    -28247, -28783, -30078, -32221, -29496, -29990, -28559, -26550, -23771, 
    -19447, -16358, -13326, -9404, -5069, -1678, 4432, 8132, 11612, 16386, 
    19644, 22045, 25720, 27404, 29787, 29794, 30594, 31407, 29353, 28251, 
    26277, 22780, 20630, 17342, 13095, 9716, 5590, 300, -2629, -6631, -12002, 
    -17451, -19710, -23198, -25634, -28522, -28880, -30639, -31501, -30086, 
    -29101, -28690, -26379, -24574, -20399, -16003, -12874, -10275, -6001, 
    -895, 3538, 7190, 11831, 15529, 19814, 23100, 26427, 27173, 28847, 29973, 
    30705, 31634, 29959, 28771, 26161, 24328, 20729, 17517, 15005, 10672, 
    4947, 1751, -3306, -8429, -12554, -15774, -19415, -23231, -24421, -27076, 
    -29480, -31690, -29683, -30794, -29643, -27127, -27215, -24663, -21998, 
    -18703, -12800, -9251, -6557, -890, 2957, 6864, 11728, 15283, 19793, 
    23569, 25843, 27432, 30159, 28550, 31180, 31561, 30161, 28428, 27270, 
    24461, 19705, 18446, 14321, 8638, 7051, 1221, -1996, -8100, -11380, 
    -15296, -20676, -22104, -25728, -28728, -29231, -30503, -30807, -30334, 
    -28768, -28116, -24950, -24228, -22019, -17747, -14368, -11196, -6753, 
    -2506, 2426, 8503, 11800, 14495, 19445, 22950, 24310, 26676, 29401, 
    31141, 32046, 29762, 29311, 27972, 27702, 24708, 21141, 19136, 13822, 
    9509, 7165, 1512, -3533, -7090, -10298, -15045, -18621, -22331, -24476, 
    -25886, -28780, -29738, -30120, -30819, -29904, -29163, -27707, -23706, 
    -21479, -19133, -13730, -10797, -7318, -359, 2298, 8309, 9976, 15306, 
    18134, 21167, 23130, 27153, 29886, 29444, 29538, 30505, 30367, 28566, 
    26222, 24015, 21891, 19227, 15143, 9779, 6313, 1912, -2624, -6062, 
    -10835, -14427, -18543, -21771, -25156, -26171, -28640, -29837, -31117, 
    -29908, -30399, -30431, -27705, -25174, -23477, -19388, -16041, -10948, 
    -6090, -2939, 1568, 4708, 9627, 15205, 19064, 22539, 25242, 25485, 29880, 
    30949, 30868, 30946, 29647, 28921, 27835, 23919, 23686, 18575, 15072, 
    11919, 5891, 4103, -2592, -4566, -11370, -14602, -19205, -20591, -24879, 
    -26092, -27530, -29687, -30041, -30930, -31047, -29081, -28020, -26437, 
    -20850, -18853, -15105, -10529, -8519, -2632, 1196, 5227, 9528, 14156, 
    17568, 21760, 23764, 28038, 28869, 29872, 29645, 31176, 31360, 29766, 
    27441, 25472, 22901, 20245, 16930, 10126, 7626, 2024, 353, -5106, -10575, 
    -12578, -16011, -20949, -24094, -26049, -28980, -29693, -31963, -32122, 
    -30546, -27693, -27092, -27265, -23179, -19910, -16261, -12108, -7541, 
    -2627, 1176, 5681, 10873, 13458, 18064, 20506, 23087, 26947, 29468, 
    30050, 31334, 30148, 30552, 30022, 28024, 25670, 23124, 19409, 16188, 
    10558, 7210, 4303, -649, -4061, -9406, -13288, -16385, -21332, -22273, 
    -26357, -28989, -29519, -30423, -29959, -30156, -29585, -27027, -26407, 
    -24037, -19846, -16986, -12623, -8644, -3479, -984, 3839, 10179, 14121, 
    17498, 20207, 24480, 26186, 29098, 28520, 31602, 30879, 30547, 28352, 
    27238, 26996, 23943, 20922, 14755, 12223, 8829, 5662, 1370, -4504, -7748, 
    -12989, -16721, -21098, -21839, -25714, -27486, -30195, -30307, -30731, 
    -31082, -28767, -26842, -24917, -23148, -19787, -17142, -12064, -8783, 
    -3748, -584, 2918, 7262, 12799, 17435, 20196, 24852, 24396, 28704, 29663, 
    31073, 29575, 30772, 30013, 26842, 25124, 24798, 19466, 17291, 14572, 
    8121, 4491, 688, -4207, -9317, -12302, -16771, -19662, -22868, -25989, 
    -28619, -30890, -30400, -31524, -30375, -29541, -29786, -26074, -23754, 
    -20478, -18068, -12910, -8817, -3094, -1811, 4850, 6888, 10881, 16255, 
    19229, 22759, 24444, 27354, 29748, 32139, 31507, 31550, 29961, 28030, 
    25254, 24424, 20039, 17313, 14921, 9607, 6322, 475, -3582, -7617, -12256, 
    -17009, -20076, -22163, -25825, -27927, -28099, -29761, -30831, -30946, 
    -29675, -29802, -26074, -24654, -22454, -18226, -14206, -8931, -5840, 
    -1272, 3064, 8281, 11382, 16372, 18480, 22020, 24983, 26088, 30121, 
    29433, 31403, 30666, 30384, 28229, 24948, 23747, 21029, 17799, 13135, 
    10624, 5440, 820, -2455, -7368, -10810, -14556, -19469, -22529, -24452, 
    -29144, -28937, -30661, -31873, -30686, -31246, -29536, -26595, -24361, 
    -20858, -19094, -13941, -10385, -5589, -1148, 3953, 5812, 11502, 15472, 
    18220, 21211, 25149, 27378, 30473, 30921, 32234, 31092, 28656, 29083, 
    27563, 24372, 20105, 18269, 13888, 10025, 4881, 1872, -3145, -7532, 
    -11512, -15129, -19418, -23106, -25986, -26516, -27975, -30396, -30868, 
    -31484, -28669, -29697, -26448, -23844, -20199, -17927, -13813, -9983, 
    -7263, -1470, 3128, 6679, 10238, 14700, 17891, 22130, 24883, 28281, 
    27466, 29917, 30473, 30733, 30034, 28373, 26062, 24639, 21604, 18857, 
    12889, 10550, 4843, 616, -2371, -6236, -11292, -16310, -19327, -21841, 
    -24774, -26464, -29283, -31023, -31046, -31268, -30236, -28614, -27346, 
    -23877, -22351, -18477, -14786, -10545, -6856, -649, 2024, 7305, 9654, 
    14743, 17639, 22223, 22818, 28664, 28414, 29094, 30011, 31138, 30730, 
    28972, 27116, 24942, 22009, 18102, 15675, 11027, 6176, 795, -1134, -6147, 
    -10097, -12714, -18029, -20382, -24265, -26983, -30059, -30198, -29934, 
    -32071, -29623, -30061, -28473, -24858, -22846, -16960, -15073, -10524, 
    -6663, -2332, 684, 6156, 9879, 15298, 17413, 22055, 23399, 27263, 29488, 
    30952, 30339, 30156, 29650, 29801, 28133, 24750, 22186, 19925, 15083, 
    11647, 7523, 2909, -1483, -4814, -9352, -15210, -17861, -21717, -25284, 
    -26665, -28108, -29944, -30467, -31069, -30345, -30178, -29321, -25153, 
    -23192, -19586, -14426, -11568, -7681, -3285, 1722, 4442, 9410, 14047, 
    17535, 20669, 24082, 25038, 28430, 29771, 29772, 29672, 29926, 29927, 
    26781, 25001, 23565, 18782, 14896, 12970, 7844, 1490, -1832, -4897, 
    -10920, -12347, -17522, -20485, -24478, -26466, -29765, -30403, -31174, 
    -29635, -29892, -28210, -29144, -25746, -22282, -19773, -15041, -12995, 
    -8309, -3170, 198, 4361, 8835, 12936, 16831, 22089, 23432, 26100, 28999, 
    28311, 30147, 31181, 30246, 28261, 28126, 24170, 23851, 19279, 16074, 
    12460, 8422, 3277, -517, -5490, -8765, -13885, -17123, -20998, -23011, 
    -26086, -27230, -29865, -30501, -31187, -31555, -28010, -28808, -25678, 
    -23853, -20541, -15162, -12549, -7436, -5078, 2148, 4915, 10187, 14239, 
    16105, 19962, 22897, 24553, 27440, 30742, 31309, 30892, 31244, 30566, 
    27934, 25503, 23888, 20352, 16091, 14170, 8580, 4097, -1798, -3607, 
    -8301, -13187, -15904, -20776, -22093, -24758, -26917, -29193, -31571, 
    -31764, -31479, -30312, -29271, -25738, -23058, -20468, -16772, -13501, 
    -8006, -4860, -100, 3096, 8023, 14189, 17238, 20607, 22266, 25812, 27632, 
    29212, 30946, 31824, 29756, 30698, 28548, 26292, 24355, 20311, 17525, 
    12653, 8649, 4115, 973, -3954, -9332, -14221, -16296, -19826, -22916, 
    -24445, -27760, -28955, -29973, -30518, -29514, -31305, -26635, -24860, 
    -22650, -21508, -16298, -12797, -7468, -6277, -668, 4280, 9184, 13639, 
    15993, 18912, 22416, 26657, 28519, 28847, 29758, 32100, 30053, 30250, 
    28997, 26087, 23877, 21421, 16709, 13328, 8616, 5131, 917, -3906, -8865, 
    -12423, -14860, -18727, -21236, -25761, -27211, -28978, -29237, -30969, 
    -30844, -29503, -29089, -26725, -24420, -19809, -17156, -14930, -10097, 
    -5457, -1895, 4921, 9300, 12654, 15675, 18441, 21754, 25860, 26627, 
    29474, 30338, 30246, 31303, 28535, 28226, 26643, 24459, 20372, 17171, 
    13489, 8171, 5417, 1227, -2305, -8347, -12966, -15081, -19180, -23808, 
    -24359, -27705, -28399, -31513, -31097, -30603, -31123, -29614, -25484, 
    -23037, -20323, -17536, -13304, -8682, -5049, -1637, 3947, 7688, 10475, 
    15076, 18049, 21866, 24631, 27788, 30187, 29696, 30006, 32007, 31531, 
    27861, 27509, 24755, 21595, 17324, 13911, 10209, 7697, 1430, -2903, 
    -7737, -10628, -15393, -19181, -22560, -25330, -26169, -30079, -30706, 
    -29453, -30072, -28747, -27780, -26926, -23712, -20839, -18101, -14796, 
    -9491, -7479, -2421, 3910, 8163, 10817, 15341, 19353, 22987, 24633, 
    27304, 29556, 30760, 29123, 32021, 31192, 28622, 26958, 24514, 20953, 
    17088, 14437, 10200, 7195, 613, -2745, -5933, -10989, -15169, -18427, 
    -21736, -25013, -27284, -28021, -31346, -29829, -30057, -29077, -28688, 
    -25456, -25355, -21721, -18498, -14309, -9102, -6707, -1649, 1952, 5737, 
    11134, 14709, 18180, 20921, 25503, 28485, 29214, 30069, 30947, 30211, 
    28957, 28224, 28243, 24669, 21958, 20172, 14905, 10366, 6411, 2102, 
    -2425, -5544, -11266, -13439, -18343, -22740, -24405, -28111, -28298, 
    -29072, -30849, -30554, -30616, -28813, -26241, -25602, -20628, -18276, 
    -14483, -12554, -7727, -3680, 1687, 7849, 8885, 14417, 18873, 22891, 
    23833, 27663, 29210, 30230, 30307, 31316, 29645, 28489, 27908, 24964, 
    22369, 20281, 15589, 11965, 8030, 4083, -1260, -6502, -10826, -15851, 
    -16800, -21168, -23627, -26516, -27741, -28535, -31614, -30931, -29067, 
    -29531, -27032, -26331, -21301, -18239, -16757, -11162, -7660, -3216, 
    1214, 6483, 9270, 14394, 16970, 20185, 23328, 25928, 28673, 28578, 29983, 
    30973, 30953, 28389, 26904, 26958, 21675, 17976, 15206, 11021, 9281, 
    3309, -750, -4045, -10486, -14925, -18833, -19829, -24632, -26206, 
    -28045, -28753, -31972, -30564, -30977, -29747, -27696, -26051, -23395, 
    -18453, -16804, -11354, -8433, -4191, 149, 6206, 11090, 12379, 16439, 
    20532, 23107, 26766, 27971, 30615, 29478, 31339, 31910, 30183, 27636, 
    24870, 24215, 19516, 16217, 11010, 7492, 4169, -730, -4667, -10381, 
    -13542, -16782, -20905, -22752, -26674, -27098, -30315, -29426, -31937, 
    -30953, -28745, -26609, -24436, -22540, -18639, -17927, -13451, -8562, 
    -4144, 294, 5030, 7674, 12253, 17210, 19750, 22991, 27410, 28412, 29925, 
    30815, 30964, 29199, 29542, 28566, 27022, 22361, 21643, 17982, 11774, 
    9027, 3939, 98, -5646, -10249, -11982, -15592, -20533, -23988, -25328, 
    -28234, -29475, -30094, -30596, -30169, -29511, -27264, -25424, -22521, 
    -19077, -15806, -12331, -7081, -4335, 5, 5913, 8695, 12440, 17827, 19564, 
    22496, 25209, 27582, 28402, 30228, 29721, 30466, 30435, 28066, 26294, 
    23930, 19178, 17191, 13474, 8583, 4768, -742, -4191, -8262, -12958, 
    -15858, -21361, -21986, -25908, -26696, -28290, -31036, -30860, -30088, 
    -30872, -27859, -27167, -24639, -20040, -16774, -12164, -9913, -4831, 
    -270, 2512, 7090, 13296, 15635, 19659, 23209, 25496, 27811, 28811, 30738, 
    31318, 30223, 30400, 27762, 26419, 24683, 19931, 17551, 14244, 8840, 
    3802, 668, -3196, -8119, -11581, -16782, -18372, -22126, -24078, -27639, 
    -27723, -30245, -28997, -30575, -29866, -28895, -28025, -23388, -21723, 
    -17668, -14432, -9501, -5869, -700, 3289, 7678, 12301, 16208, 18979, 
    22916, 25619, 28590, 28782, 29009, 29760, 29968, 30558, 27634, 27013, 
    25046, 20221, 17578, 15127, 10435, 6112, 975, -3884, -7184, -13021, 
    -15735, -20197, -21404, -26538, -27727, -29044, -31318, -31839, -30420, 
    -30402, -27621, -27235, -23983, -20759, -17329, -14221, -9642, -5840, 
    -1391, 2699, 6709, 10469, 15085, 20407, 22842, 25709, 28227, 29873, 
    30834, 32274, 30612, 29642, 28401, 25577, 24957, 22698, 17370, 14798, 
    9264, 6085, 691, -2814, -8441, -9819, -16081, -18428, -23783, -23997, 
    -28287, -27912, -31109, -31204, -30303, -31037, -28519, -26038, -23466, 
    -20841, -16871, -14459, -9972, -7544, -2190, 4331, 7852, 10475, 14003, 
    19436, 22749, 25357, 26957, 28657, 29225, 31191, 30233, 29151, 29527, 
    26826, 24075, 20635, 17083, 13530, 10748, 5226, 3181, -2972, -5710, 
    -12205, -14096, -17661, -21051, -24848, -27590, -30334, -31192, -29329, 
    -30409, -30735, -29031, -27357, -23372, -22432, -18510, -15409, -10394, 
    -7403, -2970, 2764, 6595, 10408, 15259, 17593, 23322, 25636, 27629, 
    28704, 30621, 29783, 29158, 30282, 28702, 28165, 25357, 22520, 18851, 
    14734, 10618, 6157, 1488, -2043, -6301, -10830, -15537, -19390, -20795, 
    -25217, -27207, -28299, -30380, -29803, -30475, -31215, -29071, -26264, 
    -23473, -20753, -19059, -14346, -10150, -8519, -2476, 1880, 5276, 10662, 
    15599, 17910, 20283, 24791, 26189, 28763, 30043, 30676, 30617, 30360, 
    28577, 28046, 24594, 21782, 18465, 14339, 12100, 8086, 1622, -2533, 
    -5536, -9993, -13822, -18049, -22406, -24202, -25248, -28370, -29374, 
    -28999, -30319, -30082, -29373, -28098, -25702, -21742, -19442, -15438, 
    -11264, -6991, -3443, 1549, 6222, 10599, 15151, 16006, 21365, 25135, 
    26931, 27919, 28555, 31547, 29300, 30440, 29458, 26031, 26617, 22373, 
    19911, 16901, 11547, 7606, 2586, -1009, -4541, -8838, -13399, -18895, 
    -22709, -24020, -25654, -28278, -30099, -29337, -30856, -29970, -30313, 
    -28250, -24965, -21569, -19158, -16799, -10823, -5926, -2707, 1375, 6369, 
    10575, 12287, 17900, 20022, 23881, 26179, 28354, 28834, 30064, 30493, 
    28825, 29234, 26272, 26078, 23042, 20257, 16251, 12721, 8731, 3130, 
    -1135, -5180, -10282, -14731, -17551, -20128, -22907, -26559, -29002, 
    -29657, -31701, -31720, -28760, -29301, -27382, -25710, -21618, -20936, 
    -15514, -11209, -8563, -5092, 32, 4976, 9585, 11591, 18459, 19184, 24880, 
    26580, 27898, 28336, 30277, 29877, 31593, 28695, 28840, 26579, 24470, 
    19331, 16454, 11448, 9128, 4141, 1, -5493, -9028, -13365, -16919, -21312, 
    -24010, -26679, -27882, -30343, -30246, -31304, -29703, -30286, -29650, 
    -25942, -22590, -20336, -17032, -11418, -9932, -4740, -43, 3109, 8250, 
    11906, 16302, 19566, 22671, 25624, 29560, 29433, 31039, 31693, 29592, 
    30504, 28354, 26314, 22294, 21134, 17317, 12810, 7231, 4708, -180, -3381, 
    -7286, -13099, -17386, -19053, -23429, -24363, -27787, -28763, -31034, 
    -31182, -30648, -30435, -27801, -26979, -22957, -21104, -17853, -12440, 
    -8452, -3877, -107, 4563, 9390, 13339, 16547, 21070, 22951, 25102, 27287, 
    29672, 31414, 31457, 31302, 29927, 27641, 26511, 22972, 21149, 16887, 
    12893, 10835, 3537, 1022, -4666, -7640, -12424, -17245, -19309, -22028, 
    -24939, -27309, -30684, -30340, -31298, -31268, -30642, -27654, -26210, 
    -23758, -21848, -15884, -13409, -8268, -6768, -1387, 2687, 8367, 12110, 
    15570, 17881, 23718, 26406, 28145, 29010, 29790, 29267, 31105, 30323, 
    29568, 27744, 24183, 20402, 19311, 13068, 10182, 3760, 480, -2493, -6430, 
    -12831, -15521, -18166, -22207, -25204, -28951, -29469, -30355, -31453, 
    -31035, -29010, -28330, -25899, -24141, -20708, -17420, -14105, -10443, 
    -4471, -1851, 3679, 8237, 12410, 16406, 20287, 21160, 23475, 27369, 
    28784, 30271, 30983, 31456, 29033, 30318, 27704, 25842, 21520, 18868, 
    14358, 10861, 5596, 2917, -3855, -7025, -12047, -15312, -18159, -23214, 
    -23682, -28367, -29689, -30136, -31378, -29617, -30351, -28249, -26891, 
    -25180, -22441, -17385, -15938, -8503, -6706, -3170, 2717, 5243, 10571, 
    14473, 19658, 22863, 24348, 27626, 30229, 31084, 31406, 29590, 29934, 
    27707, 26259, 25061, 22371, 18514, 15200, 11750, 6324, 1071, -2182, 
    -6385, -11373, -15919, -17881, -20818, -25518, -27396, -28455, -30623, 
    -29297, -29741, -30962, -27740, -26736, -24443, -22676, -16991, -15698, 
    -9739, -8128, -684, 2381, 4921, 11776, 15874, 18993, 21642, 25620, 26710, 
    28584, 30015, 30036, 30988, 30301, 29056, 28067, 24252, 22822, 18776, 
    14570, 11673, 5560, 1999, -2898, -7381, -9902, -13279, -17601, -23029, 
    -24557, -26229, -28341, -30438, -30734, -30782, -29083, -28220, -26039, 
    -24682, -21811, -18565, -15322, -12296, -7564, -1071, 1442, 6639, 11311, 
    14404, 18319, 21372, 23323, 26122, 28122, 29330, 30775, 31195, 30471, 
    29388, 27248, 25123, 23234, 17838, 16549, 11649, 8144, 2382, -2817, 
    -6331, -10882, -14442, -17627, -21600, -24758, -27672, -27476, -31874, 
    -30572, -30641, -30065, -29945, -27538, -25481, -21894, -18899, -14628, 
    -11898, -6359, -3549, 627, 5117, 10308, 12749, 17055, 21512, 23329, 
    25547, 29462, 30509, 31438, 32204, 31362, 29970, 26508, 26090, 22476, 
    18898, 16909, 12785, 9021, 2202, -1119, -4335, -9115, -13706, -17111, 
    -20371, -23242, -26425, -29540, -29896, -30592, -30030, -30613, -30223, 
    -27885, -25124, -22060, -18673, -16245, -11011, -9158, -2965, 2110, 5094, 
    9622, 14061, 17874, 20593, 24060, 24639, 28072, 30435, 30267, 31093, 
    29578, 29163, 26661, 25016, 23219, 19558, 16437, 13683, 8749, 4328, 
    -1100, -5500, -9971, -11966, -17287, -19404, -22963, -25972, -27057, 
    -30769, -32241, -31442, -30746, -27963, -27419, -24900, -22215, -18709, 
    -15440, -12926, -9605, -3089, 702, 4386, 9074, 13056, 18375, 21137, 
    23965, 26258, 27823, 28770, 30015, 31534, 29502, 30268, 29242, 25363, 
    23149, 20152, 16267, 13186, 7139, 3902, -737, -3991, -8042, -13240, 
    -17353, -19036, -24499, -26874, -27906, -30358, -29852, -30800, -30677, 
    -28696, -26799, -26111, -23326, -20642, -15714, -12455, -7646, -3156, 
    -143, 3680, 8109, 11857, 17860, 20506, 22700, 25600, 26857, 30922, 31825, 
    31470, 31597, 29448, 28957, 26317, 23179, 19953, 16627, 12638, 10003, 
    4461, 698, -4610, -9056, -13903, -16728, -20534, -24151, -25215, -27934, 
    -29848, -29667, -30990, -30131, -30645, -28029, -25612, -22366, -22222, 
    -17681, -14329, -9815, -6321, -56, 4198, 7958, 12084, 17764, 20709, 
    23742, 26084, 28228, 29192, 30574, 29749, 29926, 30398, 28909, 26005, 
    23518, 20627, 17032, 13774, 8225, 4395, 1395, -3026, -9516, -11841, 
    -17753, -19458, -24198, -25168, -26780, -28611, -30426, -30616, -30094, 
    -30737, -28179, -27411, -23292, -20885, -16182, -13177, -10574, -5220, 
    -2269, 2881, 7452, 12234, 15776, 18255, 22938, 25561, 26742, 30059, 
    29154, 30339, 30571, 29338, 30127, 26198, 23140, 21467, 17940, 14185, 
    10748, 6263, 1069, -3448, -7918, -12217, -15302, -18946, -22243, -26773, 
    -28644, -29250, -29734, -30719, -31151, -31081, -27220, -27525, -25185, 
    -21685, -19295, -14856, -9122, -4995, -1029, 2708, 8082, 12382, 16982, 
    20760, 21809, 25388, 28343, 30428, 30903, 30488, 30699, 30652, 28365, 
    26800, 24596, 21887, 18035, 13947, 9073, 6169, 2626, -3729, -8690, 
    -12312, -16017, -20162, -22442, -25858, -28017, -29491, -30919, -32271, 
    -30385, -30378, -28538, -26529, -24481, -22411, -19223, -13524, -9196, 
    -5964, -592, 3018, 6905, 10613, 15339, 18356, 22900, 25405, 26259, 28419, 
    29590, 29805, 30162, 28982, 27883, 27618, 22790, 21514, 18790, 14001, 
    11196, 6001, 1674, -2328, -7167, -10213, -15263, -19071, -21946, -24167, 
    -26961, -28189, -30917, -32219, -30398, -29450, -28297, -27064, -25467, 
    -20547, -18084, -13910, -11583, -6208, -1675, 3010, 6460, 10626, 15503, 
    18741, 20740, 24249, 25246, 29748, 30026, 31047, 30993, 31650, 29525, 
    27713, 26323, 21702, 18849, 14040, 10991, 7660, 2744, -1882, -8108, 
    -10070, -15414, -19228, -21136, -24426, -25687, -27917, -30045, -29717, 
    -31350, -29452, -30555, -25979, -25987, -22677, -19224, -15219, -11015, 
    -8555, -1974, 847, 6707, 11363, 13357, 17634, 21470, 25017, 28443, 30306, 
    29312, 30728, 32474, 30071, 29918, 28154, 25848, 20762, 19553, 15743, 
    11451, 8777, 3956, -1597, -5812, -10375, -15432, -17859, -22717, -23951, 
    -27208, -28341, -30578, -30924, -29299, -30586, -29802, -28346, -25028, 
    -21327, -18990, -16874, -11025, -6641, -3017, 1974, 6196, 9767, 12949, 
    19234, 21184, 22955, 27580, 27423, 30636, 30618, 31591, 28986, 29950, 
    28434, 26109, 22293, 20291, 15806, 12520, 7633, 2542, -1797, -5552, 
    -10178, -12630, -17689, -19602, -24286, -26948, -29776, -30005, -28980, 
    -30579, -29348, -28994, -28923, -24942, -22828, -20392, -15045, -12093, 
    -8419, -3899, -220, 6640, 8860, 13834, 17371, 20705, 23752, 25793, 28681, 
    29383, 29307, 30763, 30495, 29127, 28265, 26940, 21655, 19174, 15982, 
    12004, 9567, 3803, -1157, -4660, -8065, -14611, -15935, -22174, -23849, 
    -26142, -29478, -28358, -31174, -31686, -31823, -28909, -27140, -26394, 
    -23184, -20012, -17148, -13882, -7635, -3262, 432, 3383, 7865, 13452, 
    16943, 20422, 24424, 24938, 27213, 29857, 30790, 29530, 31223, 31115, 
    28850, 25156, 23051, 21012, 17076, 11858, 7607, 2344, -296, -3274, -7406, 
    -12835, -17101, -19939, -22698, -26302, -28118, -30195, -30167, -30738, 
    -30522, -29650, -27026, -27682, -23312, -20708, -16016, -12114, -8312, 
    -3715, 627, 4561, 7393, 12903, 17963, 20505, 22869, 24075, 27042, 28461, 
    31180, 31312, 30654, 29362, 27880, 25700, 23080, 19533, 16355, 12287, 
    9268, 5610, 19, -3890, -8519, -13035, -17121, -19485, -23929, -26095, 
    -27038, -27650, -30182, -29712, -30297, -28739, -27887, -26478, -23367, 
    -19489, -17039, -13453, -8866, -5087, -2151, 5059, 8286, 12549, 16613, 
    18663, 23038, 25278, 27124, 29453, 30197, 30251, 29265, 31112, 27602, 
    25055, 22965, 19931, 16124, 13176, 8458, 4438, 2107, -3632, -9073, 
    -11695, -15172, -20702, -23875, -24553, -27933, -28648, -30873, -31319, 
    -30062, -29427, -27166, -25948, -23405, -21177, -17180, -11958, -10057, 
    -3970, 163, 4672, 8064, 12914, 15513, 19091, 22137, 25303, 28235, 31052, 
    30525, 30589, 30059, 30371, 28837, 27254, 22790, 20110, 16271, 13072, 
    9343, 5313, 504, -4505, -8873, -11890, -14343, -18784, -22235, -24756, 
    -27184, -29267, -29204, -32510, -30225, -30063, -27643, -25816, -24510, 
    -21442, -17551, -12728, -9805, -5439, -1383, 4440, 8523, 11261, 14090, 
    19544, 22610, 26253, 27683, 30488, 30836, 30594, 29897, 29028, 28387, 
    26320, 24993, 22546, 17993, 15449, 10900, 5797, 1722, -2755, -7356, 
    -12392, -14990, -18353, -21025, -26356, -26232, -29324, -31521, -30086, 
    -30930, -31404, -29587, -27495, -24603, -21437, -18952, -15150, -10164, 
    -6088, -637, 2449, 7315, 11254, 13987, 17375, 20309, 24346, 27178, 30516, 
    29992, 29323, 29767, 30222, 27593, 27143, 23728, 22342, 19238, 13110, 
    10365, 6385, 2710, -2024, -5451, -10882, -14417, -18949, -22073, -24403, 
    -26885, -29022, -29175, -30725, -30757, -30851, -29223, -28079, -24426, 
    -21502, -17908, -14188, -9229, -6707, -2975, 841, 6523, 10759, 14287, 
    17008, 21333, 23481, 26577, 29905, 30778, 28998, 30991, 29321, 28795, 
    26942, 24889, 20046, 17479, 14875, 12089, 6328, 3796, -1740, -6004, 
    -11518, -14826, -18447, -23058, -24205, -27114, -28020, -31002, -30365, 
    -31751, -28795, -29344, -26446, -24315, -21229, -18750, -15716, -11020, 
    -6009, -1917, 2618, 5200, 10558, 14024, 19455, 21450, 23031, 26888, 
    28976, 29516, 31075, 30914, 29672, 29310, 27382, 24786, 22349, 19729, 
    15408, 12512, 6746, 1723, -1534, -6883, -9691, -14237, -17019, -21804, 
    -25596, -27041, -26951, -30210, -31019, -31332, -31591, -29035, -25981, 
    -25337, -21936, -18949, -15437, -10578, -6515, -2845, 2103, 6991, 8951, 
    14187, 19108, 20028, 24621, 26930, 28818, 30490, 29884, 29784, 30640, 
    30510, 26754, 25294, 22835, 19066, 15090, 11936, 7420, 3577, -2259, 
    -6258, -10268, -13471, -17645, -21065, -25150, -27665, -27444, -30056, 
    -30850, -32163, -29731, -29423, -28072, -25086, -21850, -20229, -15195, 
    -12613, -7304, -4471, 217, 5860, 9481, 13436, 17546, 19866, 22834, 25365, 
    30040, 28754, 31039, 31319, 30725, 30851, 27208, 25183, 23079, 19232, 
    16086, 12146, 8944, 3286, -1662, -6410, -9437, -13885, -17422, -20190, 
    -24745, -26152, -28788, -29190, -30307, -31173, -30931, -30205, -28007, 
    -25618, -23431, -20703, -16479, -11731, -8916, -4112, -190, 6339, 10695, 
    13040, 15463, 20701, 24607, 26112, 27133, 29423, 30518, 31117, 30195, 
    30076, 27918, 24559, 24091, 19903, 15985, 11648, 8540, 4297, -262, -4419, 
    -8103, -11703, -16838, -20876, -23094, -27195, -28934, -28861, -30937, 
    -30377, -29570, -30545, -28885, -24395, -23720, -21126, -16316, -12055, 
    -7083, -3425, -1432, 4407, 9003, 11585, 17731, 20029, 23435, 25789, 
    27619, 29510, 30146, 31801, 29330, 29045, 29404, 24953, 25068, 18946, 
    16502, 13986, 9001, 4835, 68, -4722, -8298, -12274, -15934, -19804, 
    -23331, -25678, -27960, -28978, -30829, -30762, -29076, -30442, -28771, 
    -27082, -24571, -19952, -17299, -12315, -10273, -4954, -1067, 4826, 8845, 
    12854, 16598, 19238, 21671, 25950, 27946, 28452, 31236, 30450, 30084, 
    29094, 29592, 26950, 23575, 20024, 16137, 14220, 9664, 4046, 916, -3013, 
    -8111, -11786, -16772, -21193, -21633, -24819, -28104, -28485, -30243, 
    -30480, -29838, -30670, -27799, -27784, -23963, -20555, -18628, -14762, 
    -9114, -5234, -1910, 4915, 7092, 11791, 15189, 19572, 23199, 25361, 
    25849, 30386, 31648, 30833, 29476, 28941, 29124, 25427, 23046, 20283, 
    17914, 14075, 10486, 3778, -12, -1694, -6857, -10540, -16690, -20698, 
    -23545, -25655, -26513, -28231, -31891, -29409, -29242, -31241, -27965, 
    -26720, -23321, -21419, -17375, -13203, -8512, -5896, -1133, 3158, 8062, 
    11104, 13633, 19512, 21719, 25442, 26358, 28416, 30085, 29878, 29994, 
    30839, 28392, 25639, 24224, 20876, 19124, 13254, 9819, 5979, 2716, -2542, 
    -6798, -13119, -15622, -20872, -21918, -24779, -26002, -30391, -30062, 
    -30276, -31920, -30352, -27592, -26979, -23685, -20459, -18010, -12579, 
    -9727, -5825, -1255, 3391, 6959, 12115, 16050, 17549, 21606, 25479, 
    27920, 29230, 29963, 30858, 30072, 30690, 29925, 27774, 23912, 21452, 
    18086, 13898, 11405, 5737, 2320, -1739, -7623, -9612, -16155, -17983, 
    -21971, -24218, -26819, -28678, -31310, -30581, -31342, -29656, -27931, 
    -27883, -24294, -21723, -19076, -14093, -12350, -7383, -2165, 2978, 7804, 
    10938, 13744, 18307, 21334, 25127, 27449, 28650, 29142, 30851, 29636, 
    29060, 28622, 26516, 24877, 21930, 20415, 14823, 9515, 5196, 2084, -998, 
    -5262, -11727, -14334, -18445, -22155, -24315, -26703, -30131, -30940, 
    -32467, -30741, -30301, -28593, -26622, -25548, -23184, -17855, -14391, 
    -10950, -7601, -3366, 1883, 5892, 11680, 14560, 18802, 21689, 24483, 
    26840, 29429, 30581, 31002, 31267, 30033, 28710, 27664, 25848, 21845, 
    19538, 15014, 12460, 7559, 4156, -1645, -4819, -9727, -14288, -16894, 
    -20751, -24876, -27230, -28805, -28832, -31720, -31506, -29454, -29289, 
    -28126, -26620, -22496, -19400, -16910, -11643, -7335, -2778, -424, 6703, 
    9996, 15380, 17473, 21846, 23682, 27336, 29432, 29170, 30781, 31175, 
    29871, 29133, 27296, 24630, 21156, 19503, 14643, 11223, 6718, 3656, 
    -1147, -6764, -9511, -14189, -17466, -21020, -22895, -27081, -28521, 
    -30234, -30562, -31768, -30904, -30129, -28232, -25510, -23222, -18854, 
    -16494, -12224, -7296, -3860, 1185, 5448, 9199, 13010, 16964, 20782, 
    23943, 27299, 28749, 29178, 29505, 31044, 30450, 29809, 27405, 26563, 
    22513, 20324, 15667, 11702, 7497, 3703, 168, -5279, -9953, -12121, 
    -16746, -21282, -24388, -25461, -27259, -29518, -29568, -31302, -28966, 
    -30445, -26492, -25396, -24079, -21156, -15600, -11907, -8463, -3735, 
    -146, 4994, 8675, 12645, 16637, 20130, 24243, 25319, 28567, 30111, 31283, 
    29989, 30836, 29654, 27714, 25279, 23296, 20401, 16041, 12094, 8481, 
    2731, -326, -4582, -9864, -12445, -18245, -19102, -23664, -26057, -29207, 
    -29418, -31710, -31092, -29783, -30058, -27784, -25946, -24207, -20461, 
    -15707, -11881, -9091, -5138, 1330, 4169, 7362, 12500, 16316, 20749, 
    23335, 26726, 29534, 29587, 30028, 29596, 30034, 29926, 28662, 25740, 
    22767, 20335, 17102, 12795, 7669, 4650, 275, -4639, -9628, -11270, 
    -16295, -19831, -21963, -25889, -28187, -27722, -31357, -31427, -30343, 
    -29064, -26936, -24810, -23084, -18872, -17017, -14373, -9982, -5543, 
    -482, 4998, 8675, 11321, 15627, 18782, 23225, 26304, 27711, 29609, 28961, 
    30725, 29243, 31273, 30028, 25968, 24786, 20467, 16836, 12221, 9606, 
    5199, 319, -2907, -7470, -11556, -17360, -18433, -21303, -24111, -28462, 
    -29698, -30956, -30493, -31049, -30088, -28814, -25443, -22893, -20420, 
    -16659, -12485, -8576, -6178, 116, 1962, 7480, 11475, 16734, 20676, 
    22453, 25486, 27527, 30687, 28548, 31757, 29755, 30278, 27111, 27454, 
    24555, 21797, 18214, 13829, 10630, 6957, 2377, -2397, -5949, -11506, 
    -15173, -18722, -22695, -25455, -29104, -29922, -30996, -31221, -29322, 
    -29333, -28091, -25983, -23569, -19684, -17127, -13574, -9083, -6013, 
    -922, 3836, 5699, 9928, 14965, 18842, 22473, 25748, 27025, 27413, 31431, 
    30262, 30358, 29145, 29770, 25625, 23973, 22542, 17610, 13175, 10865, 
    6658, 2172, -2740, -7259, -10919, -14955, -20042, -22921, -24732, -26362, 
    -29577, -30180, -31121, -31188, -29491, -28346, -26087, -24206, -20076, 
    -17701, -14506, -9767, -5928, -561, 2520, 8032, 10106, 14164, 17363, 
    21909, 23474, 27911, 28829, 29383, 31933, 32012, 29320, 28472, 27060, 
    25170, 21978, 17986, 13662, 12098, 7311, 2241, -1434, -5139, -10270, 
    -15365, -18060, -21500, -24848, -28156, -28964, -29959, -30117, -30309, 
    -29842, -28641, -26496, -22952, -21474, -18006, -14343, -12109, -7547, 
    -1471, 1686, 5501, 9928, 14403, 18339, 21970, 23747, 27603, 27774, 30601, 
    31832, 30417, 28536, 27904, 27325, 23534, 21844, 18295, 14602, 11304, 
    6479, 3764, -1427, -6420, -12211, -14249, -17657, -20362, -24222, -26305, 
    -28272, -29847, -31063, -30255, -30419, -29996, -27147, -25217, -21979, 
    -18195, -13900, -11006, -8661, -2002, 2145, 5159, 10773, 14718, 17477, 
    21668, 24510, 26357, 28037, 30134, 30142, 29435, 30982, 27611, 27219, 
    25516, 23391, 17912, 14319, 11157, 7414, 1782, -1689, -6410, -9959, 
    -12941, -17209, -20141, -24119, -25603, -28850, -30978, -31054, -30338, 
    -30849, -28759, -27678, -25123, -22098, -19581, -15785, -12679, -6932, 
    -2172, 336, 4918, 10369, 13421, 18605, 20323, 25518, 28071, 28292, 30372, 
    29936, 30725, 31693, 29362, 27125, 25143, 21989, 18668, 14720, 12592, 
    8318, 3238, -1869, -5584, -9198, -13272, -18577, -22757, -24812, -26742, 
    -29106, -30455, -30693, -31371, -31605, -29885, -28474, -26318, -23555, 
    -19967, -15221, -12249, -7942, -4327, -41, 4791, 8836, 13777, 16647, 
    21535, 23188, 25055, 26896, 29942, 30559, 32602, 29633, 28475, 28677, 
    24752, 22624, 20538, 15668, 12677, 8619, 3741, 322, -5371, -9671, -13117, 
    -16232, -20903, -24159, -27203, -28702, -29770, -30264, -32188, -29924, 
    -29623, -26325, -26358, -22794, -19140, -16612, -12597, -8476, -2621, 
    -233, 5988, 8384, 13634, 16985, 21090, 24400, 25076, 28170, 29622, 30273, 
    30357, 30562, 29930, 28145, 26058, 21882, 20768, 16626, 13694, 8925, 
    4644, -393, -6390, -8616, -12158, -15996, -21048, -22516, -26529, -27362, 
    -30113, -30244, -30535, -29816, -29764, -28081, -26833, -22441, -19054, 
    -15596, -12643, -9455, -4058, -1612, 3717, 8663, 13984, 17454, 19696, 
    22884, 27376, 28745, 29974, 30330, 29700, 31927, 29013, 28796, 24669, 
    24420, 20240, 15896, 12265, 8541, 4373, 326, -3257, -8599, -12283, 
    -17360, -20279, -24240, -26243, -28099, -30114, -30394, -30293, -31168, 
    -31005, -27853, -24550, -21864, -20579, -16609, -13578, -7950, -3424, 
    592, 2806, 7441, 11530, 17040, 19643, 23717, 25427, 28693, 30467, 30797, 
    30546, 30596, 30334, 27464, 25443, 22028, 19681, 17122, 15236, 8354, 
    4828, 139, -3229, -8313, -12659, -15713, -18613, -24132, -26382, -27287, 
    -27944, -31256, -31676, -31022, -28746, -27475, -26505, -23793, -20764, 
    -17837, -13927, -9145, -5283, -243, 3672, 8573, 12103, 16310, 20989, 
    22619, 24742, 28568, 28082, 29784, 29774, 30089, 31393, 27883, 26304, 
    24680, 21188, 17830, 14231, 9310, 5611, 402, -2552, -7494, -11115, 
    -16723, -20144, -23506, -24432, -26608, -29750, -30307, -31644, -31133, 
    -30756, -28288, -26501, -23900, -20290, -18090, -14825, -9610, -5711, 
    -1290, 3395, 8116, 10593, 15433, 19216, 23651, 25209, 27896, 29046, 
    29963, 31259, 31804, 28958, 28246, 26801, 25021, 21505, 16919, 14163, 
    10447, 5580, 547, -2189, -6476, -11831, -14276, -19106, -21501, -24501, 
    -26060, -29417, -30271, -30626, -30492, -30601, -27292, -26927, -24232, 
    -21694, -16347, -16049, -10225, -5564, -2943, 4035, 7152, 11177, 15591, 
    19877, 21433, 24333, 29027, 28999, 30977, 30162, 31549, 28875, 29661, 
    26511, 24554, 22299, 17761, 14591, 12230, 5823, 1673, -2625, -6234, 
    -12152, -15538, -19493, -22406, -25575, -27160, -29618, -30417, -30019, 
    -29990, -30176, -29349, -26052, -23757, -20298, -19580, -14485, -10155, 
    -4820, -2550, 2996, 6642, 10149, 14071, 19724, 21745, 23867, 28813, 
    29584, 31111, 29762, 29237, 30096, 28580, 26789, 24369, 22461, 17239, 
    13941, 11662, 6347, 1894, -3081, -5035, -11254, -14042, -18203, -22106, 
    -23865, -26914, -28383, -30004, -30170, -31724, -29662, -28753, -27181, 
    -24980, -22847, -19966, -14747, -11024, -7119, -2236, 2334, 5678, 11302, 
    14426, 18447, 20827, 24303, 27332, 27344, 30396, 30605, 32220, 29619, 
    28165, 26248, 25090, 21593, 17591, 15153, 12431, 8080, 2849, -3122, 
    -7225, -11531, -15720, -17852, -22218, -23437, -27818, -29474, -28324, 
    -30784, -29101, -29633, -28238, -26918, -25490, -21930, -17274, -14999, 
    -11853, -7299, -3598, 2029, 7035, 9726, 14763, 18253, 21137, 24699, 
    26362, 29353, 29349, 28871, 30966, 30835, 27797, 27377, 24408, 22985, 
    20301, 15324, 11268, 8595, 4066, -892, -5293, -8789, -12964, -16722, 
    -21387, -23970, -25040, -27963, -31075, -31809, -30424, -29772, -29290, 
    -27238, -25529, -23336, -18440, -16607, -10334, -8566, -2895, 549, 4724, 
    10103, 13053, 17161, 21341, 23980, 27407, 27535, 29170, 29826, 30587, 
    29976, 29595, 27156, 25779, 24468, 19485, 16225, 12960, 7029, 4616, 
    -1539, -5194, -10165, -13574, -16722, -20675, -24579, -27099, -29364, 
    -29987, -29009, -30534, -30009, -28810, -28602, -24396, -23401, -20099, 
    -14832, -12333, -9051, -4215, 752, 4115, 7595, 11933, 17314, 21360, 
    23674, 27271, 26921, 29516, 31602, 31362, 29327, 30835, 28543, 27195, 
    24321, 20078, 16845, 11842, 8538, 4292, -857, -5490, -7797, -11898, 
    -16246, -19730, -24223, -26537, -28402, -29594, -29418, -31500, -30197, 
    -29837, -27469, -25110, -23750, -18859, -15260, -12754, -8309, -3963, 
    -225, 4641, 7108, 11376, 15357, 21119, 24356, 24813, 28726, 29664, 29912, 
    30141, 30497, 29487, 28168, 26985, 24744, 20530, 17111, 13612, 10765, 
    4275, 1420, -4208, -9370, -12921, -15214, -19251, -24538, -25446, -27178, 
    -29800, -30377, -30750, -30287, -29442, -29800, -25949, -23202, -22016, 
    -15768, -13811, -8442, -5008, -236, 3408, 9038, 12536, 15617, 20744, 
    23526, 25285, 26527, 29191, 30004, 31009, 31087, 29289, 28785, 25213, 
    23187, 22238, 17237, 13913, 9269, 5412, 1469, -4214, -8881, -12155, 
    -16690, -20065, -23462, -26553, -26576, -28330, -30153, -29152, -30972, 
    -30446, -28165, -28031, -23761, -19915, -18094, -12660, -9898, -6035, 
    -1246, 4111, 8128, 11380, 17554, 20268, 22741, 24727, 27243, 30130, 
    30972, 32091, 30608, 28747, 29882, 26553, 24578, 20998, 16585, 13349, 
    10219, 5959, 419, -1618, -8433, -12934, -15393, -18795, -22906, -24735, 
    -27894, -29547, -31252, -29830, -30946, -30294, -27898, -25881, -23507, 
    -20973, -18537, -12897, -9703, -4986, -1495, 2204, 7396, 11281, 14382, 
    18862, 22577, 24989, 26907, 28891, 30907, 31367, 30059, 31063, 27520, 
    25176, 23910, 21289, 17873, 14518, 9595, 4709, 3222, -1841, -7464, 
    -11144, -15834, -19575, -21417, -24340, -27176, -28444, -30641, -31652, 
    -30467, -29826, -27103, -25701, -23555, -21121, -16628, -15095, -9874, 
    -6892, -1740, 2559, 6302, 11794, 14510, 19403, 21021, 24941, 26783, 
    29097, 29671, 30006, 31034, 30240, 29213, 28044, 25249, 22875, 19222, 
    14683, 10736, 7500, 3429, -3143, -8017, -11554, -15964, -19035, -22831, 
    -25847, -27534, -28193, -29860, -30987, -31527, -30911, -28230, -27192, 
    -25799, -22305, -18443, -13713, -10795, -4956, -2260, 1702, 7873, 10556, 
    13942, 17007, 23003, 24798, 27605, 28667, 29198, 31363, 30464, 29740, 
    27538, 27143, 23371, 22452, 19354, 15445, 12292, 6037, 2448, -2016, 
    -6898, -11586, -14639, -18956, -22108, -24715, -26675, -27066, -30099, 
    -31694, -30733, -30658, -28778, -27245, -25302, -20391, -19056, -15840, 
    -10889, -6845, -2305, 645, 5904, 8581, 14799, 18189, 22264, 24126, 27234, 
    29725, 29445, 29755, 30394, 29570, 29595, 27644, 23740, 22594, 20321, 
    14437, 11189, 6757, 3076, -993, -5788, -10829, -13721, -18095, -20817, 
    -24294, -26294, -29177, -29684, -30367, -30159, -29716, -29963, -28000, 
    -24554, -22698, -20419, -15737, -12624, -7035, -3886, 1669, 4704, 9247, 
    14228, 16742, 19645, 25206, 27527, 28597, 29686, 31783, 29815, 30353, 
    27699, 26944, 25098, 22715, 20062, 15962, 10988, 6724, 2514, 517, -6323, 
    -9387, -14843, -18022, -21695, -23972, -26434, -28478, -29844, -29241, 
    -31194, -31354, -28371, -25966, -26837, -21326, -20616, -16492, -11504, 
    -8245, -2486, 761, 3395, 10961, 12255, 17772, 19532, 24244, 27121, 28639, 
    31257, 30546, 29580, 29167, 29812, 28239, 24892, 23163, 18059, 15895, 
    12229, 7926, 2409, -597, -5638, -8654, -14729, -17849, -19844, -23344, 
    -28051, -28262, -29273, -32117, -30831, -29357, -29506, -28826, -24245, 
    -21371, -21057, -17209, -12742, -8343, -5444, 921, 4963, 9057, 13313, 
    18435, 19948, 23459, 25412, 27321, 28156, 31836, 31045, 30422, 31201, 
    28325, 26138, 22972, 20522, 15235, 12031, 7756, 4801, 943, -4069, -8684, 
    -14576, -17175, -19654, -22995, -26404, -28066, -30868, -29092, -30086, 
    -31396, -30695, -28029, -25061, -23009, -20589, -16191, -13469, -9166, 
    -4175, -268, 5407, 8866, 11738, 17378, 19702, 23279, 26015, 28077, 28261, 
    31248, 30294, 30997, 30306, 26299, 26340, 24939, 19809, 15685, 12899, 
    8427, 3696, 1264, -3612, -8000, -12461, -15650, -19171, -23810, -24325, 
    -28596, -29511, -30390, -31257, -30401, -29758, -28231, -27200, -23470, 
    -21725, -16593, -14557, -8280, -5203, -243, 3780, 7217, 11778, 15915, 
    21112, 23745, 26161, 28360, 29342, 29677, 29405, 30161, 30511, 27892, 
    27267, 22683, 20012, 16698, 13584, 10387, 5305, 431, -2995, -7761, 
    -11756, -16912, -20239, -22889, -26569, -27387, -29466, -30679, -31766, 
    -30851, -30277, -28636, -27118, -23410, -21824, -16975, -13483, -10703, 
    -5293, -983, 3956, 8408, 12109, 14802, 18682, 23493, 25032, 28592, 29603, 
    30866, 31653, 31218, 29783, 27915, 26782, 22232, 21244, 17861, 13043, 
    9099, 6987, -539, -2948, -6718, -10627, -15508, -19668, -23563, -26844, 
    -28568, -29263, -30258, -32108, -30838, -29872, -28148, -27277, -24033, 
    -22248, -17918, -15210, -9992, -5960, -1512, 4267, 8631, 11265, 16399, 
    18352, 22137, 25771, 27003, 29924, 30644, 30426, 31027, 29239, 29193, 
    25703, 24244, 20924, 18842, 13905, 10798, 4850, 2723, -4176, -8285, 
    -11399, -15406, -20333, -20606, -24521, -25911, -28406, -31464, -30665, 
    -29885, -30309, -29046, -26585, -24719, -20518, -19396, -14352, -10645, 
    -5132, -2573, 2190, 7093, 10619, 14655, 19380, 22178, 25367, 27612, 
    27877, 29045, 30665, 30384, 29586, 27905, 26446, 25168, 20424, 18859, 
    13812, 10810, 6707, 2352, -1950, -6761, -11036, -15948, -17502, -20946, 
    -24291, -27154, -28768, -31664, -30685, -31425, -30633, -29518, -26881, 
    -25002, -22372, -18628, -14790, -10161, -6788, -2052, 2448, 6938, 9121, 
    15710, 17055, 22628, 25417, 26330, 28728, 30257, 30976, 30362, 30950, 
    29607, 27246, 23764, 21489, 19560, 15696, 12230, 7617, 1014, -2536, 
    -7034, -11495, -13840, -18675, -20125, -24692, -26370, -30616, -30349, 
    -30236, -32162, -30494, -28306, -26309, -25105, -21291, -18154, -14781, 
    -10761, -5821, -2559, 1284, 5975, 11152, 13319, 16655, 21884, 24906, 
    25737, 28753, 30429, 30499, 31987, 30283, 29727, 25652, 25184, 22183, 
    19621, 16196, 11044, 7687, 3143, -1265, -5935, -11159, -13404, -17269, 
    -20103, -24580, -25369, -29149, -30882, -30162, -29388, -30066, -27919, 
    -26753, -25018, -23207, -18818, -15854, -10186, -8371, -1987, 1360, 4411, 
    10557, 14308, 17706, 20119, 24177, 26045, 29161, 30261, 29472, 29665, 
    29943, 28600, 27336, 25139, 24021, 20540, 16896, 11879, 8032, 3703, 48, 
    -5144, -8388, -13982, -17325, -20296, -24269, -26483, -27036, -29125, 
    -30823, -30759, -30455, -28599, -28196, -25989, -23095, -21046, -14737, 
    -12442, -7942, -4022, 908, 6252, 11129, 13022, 17233, 19226, 24525, 
    27237, 30094, 29604, 29307, 31281, 30231, 30435, 29175, 24673, 23050, 
    20267, 15678, 12167, 8162, 3693, -1458, -5177, -7534, -13394, -15943, 
    -20785, -23274, -25783, -28047, -29756, -29375, -29563, -30720, -28616, 
    -27421, -26702, -22877, -18802, -15168, -13753, -8645, -3843, -130, 6637, 
    7743, 13886, 16383, 20349, 25344, 24904, 28032, 29377, 30238, 31191, 
    31171, 28215, 27084, 25009, 21820, 19966, 16976, 13034, 8747, 5731, -892, 
    -5664, -7924, -11867, -17290, -20185, -22417, -26265, -27231, -30047, 
    -31095, -30992, -29244, -30870, -26917, -25732, -22609, -19324, -16894, 
    -14259, -10057, -5413, -266, 3922, 7803, 12624, 16865, 20924, 22760, 
    24992, 28262, 31016, 30423, 31316, 31865, 30860, 29234, 25811, 23404, 
    20571, 18273, 14144, 9974, 3321, -581, -2245, -8888, -12557, -17950, 
    -19804, -22533, -26214, -28847, -29375, -30119, -30339, -31429, -30542, 
    -28733, -26464, -23790, -20572, -16820, -12735, -8127, -6237, 937, 3547, 
    7511, 13982, 14953, 18999, 23301, 27026, 27697, 29635, 30394, 32596, 
    31287, 29660, 27929, 26834, 22955, 20789, 15495, 13905, 9458, 4613, 1667, 
    -3368, -7488, -10917, -16085, -20545, -23678, -25582, -27805, -29518, 
    -29526, -30511, -30685, -28508, -28826, -26924, -25415, -22201, -18384, 
    -13420, -10153, -3943, -2158, 3874, 8469, 11971, 14428, 19024, 24059, 
    24285, 28328, 28077, 29248, 29826, 30545, 30287, 29316, 27154, 24070, 
    22404, 17688, 15010, 9337, 5144, 2430, -4835, -6483, -11748, -15238, 
    -20268, -22852, -26998, -26599, -29592, -30819, -30927, -30693, -29685, 
    -27412, -25667, -24378, -21482, -18139, -13933, -9441, -5336, -1513, 
    2959, 8516, 12446, 13790, 19662, 23449, 24901, 28780, 29082, 30063, 
    31313, 30789, 29921, 28226, 25840, 23558, 21481, 18409, 13942, 11278, 
    4808, 1490, -3690, -7179, -11743, -15034, -17484, -23896, -23668, -27462, 
    -29262, -31664, -30458, -31239, -30191, -28177, -26184, -24142, -21369, 
    -18063, -13072, -9049, -6756, -837, 2877, 5695, 10447, 14342, 18593, 
    21778, 25811, 27071, 28928, 31228, 29419, 30582, 30810, 27159, 28000, 
    24869, 20479, 19137, 13319, 10934, 6831, 2405, -2884, -6695, -11687, 
    -14012, -17482, -20640, -24687, -26946, -28537, -29942, -30885, -32030, 
    -30276, -28234, -26262, -24458, -21540, -18919, -15252, -11002, -6029, 
    -706, 1897, 7556, 11778, 14200, 18792, 21312, 25120, 26756, 28085, 30901, 
    30882, 32571, 30011, 29588, 26987, 23855, 20419, 19129, 16261, 11403, 
    8495, 2856, -2815, -5423, -11643, -14895, -19480, -21378, -24473, -26531, 
    -30006, -30231, -31105, -31162, -30234, -28009, -27269, -25177, -21617, 
    -17995, -14019, -9914, -7131, -3579, 1735, 6945, 9404, 13464, 18767, 
    21990, 24216, 27051, 29701, 30963, 30298, 30172, 30051, 28841, 26952, 
    25099, 22299, 18434, 16385, 10902, 6926, 2023, -1128, -5240, -10515, 
    -14798, -17910, -19382, -25165, -26229, -29902, -29392, -31563, -31837, 
    -30691, -28003, -28353, -24723, -22907, -18988, -16882, -10401, -7837, 
    -3761, 693, 5881, 11821, 15024, 15905, 20513, 23615, 28002, 27896, 28831, 
    29755, 30744, 31577, 29567, 26036, 26704, 22196, 18433, 16466, 13297, 
    6332, 3571, -787, -4338, -9967, -15359, -17740, -20297, -22573, -26464, 
    -29060, -29876, -31365, -30146, -31437, -29934, -26992, -24865, -22856, 
    -19061, -16199, -11944, -7308, -3124, 1882, 5919, 8760, 13221, 17126, 
    20644, 22182, 27402, 28618, 30176, 30752, 31602, 29430, 29833, 28220, 
    25953, 23361, 19986, 15517, 12872, 7272, 4544, -1121, -4190, -11090, 
    -11969, -17300, -19447, -23725, -24582, -28857, -30143, -31742, -30546, 
    -28797, -28649, -27769, -26279, -23600, -19679, -14985, -11718, -8315, 
    -3981, -426, 3854, 8311, 13120, 17941, 21603, 23633, 26949, 29178, 30049, 
    31508, 30552, 29605, 29938, 27503, 26421, 22565, 19128, 16752, 11649, 
    9043, 3228, 910, -5346, -9563, -14591, -16808, -20494, -22117, -25475, 
    -27591, -29224, -32195, -30711, -30985, -29778, -28341, -24571, -23513, 
    -20482, -16251, -11819, -8296, -4397, 39, 4421, 9425, 12342, 17953, 
    21556, 23146, 26241, 28419, 30436, 31514, 32026, 30743, 29096, 26557, 
    25192, 23187, 19778, 17591, 12911, 9620, 4559, -750, -5657, -8838, 
    -12692, -15755, -19542, -22070, -25463, -27105, -27858, -31031, -30215, 
    -29238, -30944, -27242, -26255, -22829, -19439, -16751, -13352, -8397, 
    -3702, -838, 3383, 6971, 13567, 16444, 18656, 22604, 26011, 26661, 30149, 
    31732, 29433, 30401, 29395, 27684, 24820, 24463, 20704, 16654, 14224, 
    10977, 5631, 1788, -4810, -6568, -12599, -16587, -20877, -22732, -23883, 
    -28205, -28155, -30273, -31896, -29687, -30688, -28323, -26304, -23938, 
    -19333, -16734, -12944, -9377, -4592, -1588, 5069, 7962, 11211, 17176, 
    19386, 24006, 26991, 27124, 29747, 30427, 31711, 30835, 29558, 29136, 
    27345, 25823, 21415, 16388, 13600, 10273, 5975, 423, -3529, -8755, 
    -11170, -15291, -18168, -23953, -25443, -26574, -29898, -31321, -30141, 
    -29351, -28151, -28144, -27044, -22445, -21127, -16594, -15321, -9964, 
    -6020, -1006, 4509, 6497, 12662, 15245, 19190, 22359, 24400, 27127, 
    30159, 30162, 31097, 30701, 29877, 28714, 27802, 24897, 21764, 19380, 
    15148, 10027, 5684, 902, -3254, -7431, -10783, -15750, -18933, -22936, 
    -25564, -28621, -29246, -31123, -30710, -31489, -30998, -27210, -26401, 
    -25915, -21710, -17886, -15235, -11511, -6278, -2594, 4000, 6786, 12356, 
    14509, 19568, 21439, 25265, 28251, 28873, 30704, 30649, 29852, 30830, 
    28816, 28637, 24765, 21044, 18346, 14819, 10290, 5010, 3586, -2422, 
    -7437, -11486, -15478, -18962, -21076, -25379, -26978, -29580, -30475, 
    -30270, -30336, -30826, -28061, -26097, -24528, -21818, -17045, -14890, 
    -11478, -6550, -1961, 2018, 6827, 10065, 15406, 19388, 21835, 24452, 
    28513, 27296, 29228, 30473, 31749, 29274, 29356, 26412, 23213, 22446, 
    18684, 14820, 10065, 5412, 3152, -1004, -7030, -11415, -15129, -18016, 
    -21584, -25809, -27030, -29535, -31145, -31367, -31322, -29558, -28038, 
    -26706, -24402, -22817, -19060, -14639, -11018, -7207, -3881, 1077, 6872, 
    11229, 13934, 19359, 20168, 24900, 25735, 29870, 29746, 29030, 29785, 
    29693, 27953, 27199, 24835, 23408, 17775, 14214, 12101, 8168, 1442, 
    -1645, -4249, -9624, -14893, -18558, -21756, -24105, -27282, -28994, 
    -29610, -30705, -30943, -31346, -30017, -27097, -25055, -22012, -18546, 
    -15802, -11370, -8457, -2898, -474, 5730, 9285, 13757, 18194, 21446, 
    24336, 26229, 29070, 28720, 31689, 30088, 29695, 29365, 26479, 25451, 
    22981, 18791, 16521, 11699, 6685, 2292, -1575, -5698, -9408, -13342, 
    -17149, -21277, -24443, -25481, -27794, -28766, -29254, -32114, -29145, 
    -28358, -28247, -26483, -22029, -20209, -16247, -10757, -7598, -3294, 
    383, 4368, 10290, 12542, 18049, 21771, 22888, 25811, 28812, 31298, 31630, 
    31065, 30297, 29169, 27446, 25165, 22882, 20676, 15473, 12193, 7461, 
    2030, -545, -4729, -10470, -14512, -17757, -21293, -23771, -25212, 
    -26874, -30672, -29280, -30864, -30622, -30336, -27811, -25086, -23230, 
    -20908, -16122, -11460, -8404, -4566, 237, 5134, 8450, 13108, 17789, 
    19696, 24368, 27246, 28493, 30140, 31051, 31624, 30166, 29982, 27716, 
    25410, 24161, 21274, 17179, 12773, 7813, 4725, -1482, -2878, -9304, 
    -12154, -18305, -20092, -23390, -25513, -27941, -29808, -31819, -30695, 
    -30146, -29463, -28810, -25612, -22402, -19426, -16328, -13803, -7708, 
    -4851, 982, 2725, 9769, 12668, 17432, 19354, 23476, 26107, 27927, 30380, 
    28849, 31113, 29102, 28064, 28889, 25512, 23401, 19946, 17141, 13282, 
    8101, 3928, 29, -4553, -7895, -13350, -15213, -20916, -23528, -26492, 
    -27820, -30120, -30791, -30260, -31792, -29818, -29329, -26388, -23625, 
    -20883, -17481, -12562, -9640, -4894, -318, 3828, 8559, 11066, 16305, 
    19472, 23609, 25316, 27897, 29428, 31148, 30755, 31022, 30518, 28105, 
    26511, 23953, 19715, 17565, 14671, 7916, 6677, 534, -4446, -7300, -12081, 
    -16205, -18889, -22305, -23793, -26878, -29508, -28937, -30920, -32015, 
    -30069, -28288, -26400, -24352, -20260, -17383, -13256, -9288, -4655, 
    -656, 3484, 8161, 10714, 16482, 19403, 23098, 25853, 28307, 29319, 30241, 
    30660, 30916, 29251, 28575, 26761, 23394, 21144, 16996, 13116, 9556, 
    4533, 179, -4594, -7591, -11858, -16659, -19525, -20987, -24914, -28212, 
    -28151, -30960, -29271, -30018, -29352, -29734, -27055, -23335, -21396, 
    -16805, -14015, -9865, -6292, -230, 3781, 8149, 12182, 16094, 18834, 
    22304, 26728, 27751, 29116, 29678, 30281, 30483, 30802, 30192, 26726, 
    23801, 21564, 16960, 15038, 9359, 6341, 123, -2758, -6312, -9980, -15331, 
    -18857, -21977, -25211, -27622, -29508, -29346, -31515, -30839, -29726, 
    -28188, -26629, -23238, -21491, -17936, -15063, -11216, -5943, -2388, 
    2851, 6595, 11242, 15699, 18955, 20574, 24427, 26520, 28528, 30017, 
    30318, 29932, 31289, 29346, 27498, 24049, 21588, 18371, 12756, 9918, 
    6354, 1410, -727, -7150, -11432, -14997, -19030, -21450, -23239, -27377, 
    -28223, -31503, -31409, -31426, -29444, -29465, -26869, -23991, -21342, 
    -19449, -13197, -10468, -7374, -2351, 2856, 7666, 10954, 14486, 19260, 
    22354, 25524, 27148, 27127, 29634, 30228, 30990, 29707, 28001, 26845, 
    23295, 21418, 19459, 14092, 10455, 6304, 1384, -3399, -5774, -10211, 
    -13884, -17163, -21900, -24929, -27156, -27665, -29071, -31431, -30523, 
    -30265, -29209, -26489, -24414, -22485, -19834, -16158, -10946, -6958, 
    -1742, 1920, 5432, 9974, 13737, 17739, 21496, 23776, 26738, 28923, 30855, 
    31104, 31613, 29117, 28659, 26465, 25908, 22506, 18968, 17046, 12223, 
    7807, 3250, -2774, -5297, -10044, -15064, -18040, -21872, -24934, -27118, 
    -28790, -29918, -31423, -31257, -31679, -28870, -26794, -24342, -22867, 
    -17313, -14743, -12138, -6366, -4107, 1128, 6050, 9791, 13997, 18366, 
    21976, 25366, 26243, 27007, 30095, 30284, 29965, 31479, 28861, 27075, 
    24539, 20943, 20870, 15107, 11793, 8204, 3762, -1348, -6979, -8615, 
    -13016, -16167, -21716, -23424, -27602, -27281, -28423, -31294, -30630, 
    -29487, -28802, -28089, -25260, -22714, -19979, -15643, -11802, -8226, 
    -3207, 1322, 6699, 9824, 13692, 16725, 21211, 25025, 27641, 28533, 28838, 
    31017, 29834, 30090, 30734, 26914, 25464, 23694, 19123, 15668, 11328, 
    9502, 3737, 973, -5284, -9537, -13720, -17209, -20100, -23966, -27328, 
    -28649, -28724, -30352, -30854, -30436, -29669, -28504, -25614, -23122, 
    -19469, -16467, -12451, -8402, -4784, 1360, 5129, 9797, 13096, 16226, 
    22029, 22528, 24783, 26733, 28639, 30277, 31957, 30664, 30606, 27522, 
    26797, 23527, 20839, 15192, 12829, 9334, 2544, 37, -4816, -7562, -12465, 
    -17124, -20750, -24069, -26017, -28843, -29576, -30979, -31739, -30390, 
    -30412, -29145, -24395, -23196, -19564, -18178, -12772, -10128, -4147, 
    -230, 4847, 9710, 11959, 16658, 20856, 23121, 26773, 26864, 29478, 31354, 
    30706, 31132, 29549, 27384, 27311, 23997, 20352, 16671, 11893, 8927, 
    5718, -478, -4697, -7350, -12968, -16800, -20214, -21813, -25509, -28390, 
    -29140, -31157, -31356, -29925, -28654, -28064, -25179, -23482, -20567, 
    -18589, -13146, -9478, -5046, -206, 4256, 9295, 12523, 15842, 20656, 
    21933, 26485, 28916, 29606, 30673, 31643, 30094, 29803, 28683, 25053, 
    23111, 19467, 17424, 14313, 8943, 4873, 1199, -2847, -7704, -11997, 
    -15785, -19458, -22923, -25572, -27586, -28303, -29124, -31062, -30974, 
    -31325, -28321, -27055, -24084, -21645, -17968, -13856, -10471, -4032, 
    367, 2799, 8947, 12291, 16613, 20081, 22876, 24915, 27328, 28778, 31373, 
    31679, 28958, 30713, 28018, 27142, 23738, 21945, 15857, 15258, 8686, 
    5702, 497, -2735, -7707, -13630, -16206, -18434, -23090, -26002, -26040, 
    -30603, -30462, -31281, -30075, -30776, -27100, -25788, -25179, -21734, 
    -19360, -15761, -9573, -4494, -1743, 2751, 8217, 11886, 15870, 19610, 
    22083, 23979, 27697, 29048, 31101, 29846, 31654, 30032, 29980, 27974, 
    24093, 21673, 17737, 14897, 10686, 6930, 1032, -3080, -7482, -12887, 
    -13598, -18932, -21855, -25342, -28566, -29038, -30416, -29738, -29578, 
    -29959, -28631, -27082, -24168, -20926, -19626, -15578, -11777, -5881, 
    -2508, 2711, 7718, 10754, 14465, 19459, 21956, 24637, 26082, 29267, 
    30718, 31738, 30254, 30555, 29104, 27774, 23268, 21453, 18649, 14105, 
    9224, 5975, 1456, -1675, -5575, -10979, -15403, -18185, -21453, -25901, 
    -28217, -28336, -29725, -31836, -31882, -29250, -30381, -27321, -24927, 
    -22319, -18473, -15308, -10232, -7026, -1136, 2320, 6640, 12093, 13045, 
    18902, 21393, 24550, 26703, 28798, 30853, 30157, 30929, 30707, 30255, 
    25364, 24351, 22136, 19017, 15502, 11433, 8012, 3173, -1618, -6526, 
    -9633, -13326, -18494, -20284, -23716, -26735, -28844, -29564, -30400, 
    -32172, -29266, -29179, -27834, -24278, -20780, -20218, -14610, -11081, 
    -8022, -3272, 622, 5626, 9816, 13218, 17102, 21092, 23004, 26097, 28812, 
    29910, 31904, 28862, 30229, 29612, 27978, 25389, 21006, 17249, 16256, 
    13192, 7337, 2044, -2496, -5616, -9805, -14469, -17950, -20500, -24278, 
    -26339, -28408, -28922, -30639, -31109, -30326, -29768, -28241, -26099, 
    -23277, -18507, -15346, -10173, -8680, -3303, 1724, 5265, 10004, 14334, 
    17292, 20592, 23424, 25949, 29200, 31312, 29685, 29362, 29502, 30189, 
    27515, 25417, 21327, 17969, 15918, 11478, 7133, 2909, 180, -5178, -8926, 
    -12717, -17129, -22459, -23735, -25886, -28591, -30235, -30861, -30492, 
    -30413, -30504, -28092, -26808, -23042, -18489, -14949, -13043, -9430, 
    -4093, 552, 6053, 9113, 11763, 16914, 20665, 23724, 26002, 28892, 30823, 
    31816, 31518, 30369, 27688, 26855, 26119, 21968, 20286, 17964, 12332, 
    7631, 2544, -2445, -4209, -8369, -15028, -16616, -21612, -23647, -27225, 
    -27819, -29953, -28979, -29433, -29482, -30949, -28979, -24634, -22817, 
    -18619, -17764, -12593, -6869, -2203, 1136, 5914, 8634, 12142, 18606, 
    21300, 23679, 26199, 27642, 30597, 31210, 30846, 28666, 28917, 26823, 
    25208, 24050, 19224, 17233, 13084, 7406, 3205, 65, -3996, -7775, -13764, 
    -14959, -21432, -24830, -26511, -26631, -29033, -31403, -30702, -30351, 
    -30209, -27405, -25498, -21677, -18258, -17719, -13923, -7290, -4693, 
    -554, 5005, 9821, 13157, 15472, 19261, 24029, 24445, 27306, 29407, 32174, 
    31134, 29621, 30851, 28201, 26845, 23479, 20248, 16041, 13231, 8063, 
    4343, -395, -4517, -9596, -12015, -16871, -19599, -23642, -25406, -27615, 
    -30319, -29407, -30094, -32312, -29639, -29531, -26047, -21733, -19888, 
    -16480, -13009, -9608, -3678, 699, 4234, 9873, 12019, 14722, 18711, 
    23141, 25563, 26822, 29892, 30067, 30557, 29686, 30320, 29380, 26276, 
    22443, 22210, 16485, 13188, 10682, 5462, 1209, -3273, -8571, -12468, 
    -16632, -19959, -24288, -25317, -26095, -28615, -30399, -31537, -31052, 
    -30240, -27541, -26335, -23701, -22115, -16796, -12752, -10125, -3798, 
    -2646, 3243, 9310, 11476, 16119, 19991, 22935, 24471, 28367, 29768, 
    31324, 32554, 30969, 29278, 27398, 27042, 22933, 21194, 18079, 14477, 
    9804, 4614, -222, -2383, -6964, -12599, -15007, -17744, -24422, -24012, 
    -28515, -30417, -29404, -31578, -30726, -28561, -28953, -25501, -24866, 
    -20937, -18318, -14322, -9768, -5529, -2894, 1849, 9125, 11762, 17165, 
    19581, 22625, 25823, 27456, 30040, 30177, 30974, 29879, 29930, 28234, 
    26585, 23659, 21640, 16874, 13614, 10281, 6130, 1057, -2549, -6942, 
    -11989, -15300, -20275, -20648, -24447, -26624, -29422, -31605, -29646, 
    -31245, -28644, -28127, -25691, -23401, -21201, -17748, -12788, -10100, 
    -6421, -114, 945, 5524, 9817, 15842, 19292, 21728, 24285, 25907, 29119, 
    31590, 29701, 30559, 29321, 29380, 26679, 24254, 21733, 19605, 14929, 
    10582, 6491, 3255, -1410, -7355, -10448, -15975, -19550, -22300, -26515, 
    -26538, -29160, -30623, -29060, -29665, -29208, -28772, -26767, -25071, 
    -21344, -19214, -14683, -9859, -6750, -2294, 2954, 7477, 9684, 14823, 
    19396, 20608, 25136, 26812, 30078, 30923, 30711, 30650, 30955, 29156, 
    25817, 25108, 21603, 18523, 15717, 10897, 6904, 1489, -2078, -6811, 
    -10474, -15449, -17798, -22933, -23233, -25839, -27260, -30075, -30760, 
    -31763, -30727, -28094, -27323, -25190, -21942, -17923, -13257, -9737, 
    -5900, -2692, 2072, 7177, 9107, 15474, 19099, 22506, 23578, 27084, 27964, 
    30036, 29407, 29842, 30669, 27750, 26729, 24770, 23294, 20115, 16137, 
    12951, 7918, 3402, -801, -5303, -10505, -13467, -18538, -22853, -24578, 
    -28067, -27387, -30619, -31418, -31077, -31352, -28607, -28124, -24100, 
    -23085, -19269, -14765, -11816, -7041, -4278, 1207, 6333, 10910, 13312, 
    18405, 21469, 24360, 26996, 27735, 29595, 30847, 30215, 31154, 29735, 
    25866, 24639, 22447, 20911, 16992, 11599, 7433, 3505, -378, -4371, 
    -10305, -12976, -18122, -19069, -23534, -26617, -28361, -31096, -29781, 
    -31171, -31082, -31027, -26334, -23679, -22239, -19571, -14701, -11721, 
    -6719, -3875, 1261, 5091, 10547, 14357, 17608, 20892, 22062, 25655, 
    26718, 28662, 30507, 30228, 30737, 28584, 27703, 25408, 22834, 19677, 
    17005, 13102, 7947, 5579, -710, -5818, -9066, -12756, -17197, -19068, 
    -24793, -26039, -27367, -28204, -29655, -31479, -30604, -29571, -27701, 
    -26305, -22295, -18379, -17282, -12632, -8266, -3997, 1570, 4030, 10399, 
    14080, 18209, 20455, 21696, 25688, 29632, 29633, 29552, 29904, 29163, 
    29592, 27433, 24927, 23201, 21410, 17387, 12148, 7758, 3819, -1539, 
    -5076, -9825, -12202, -17106, -20095, -23425, -24954, -27515, -30280, 
    -29725, -31102, -30598, -29135, -28141, -24570, -24586, -21570, -16543, 
    -12577, -8483, -3759, -146, 3772, 8307, 12768, 15579, 20120, 23846, 
    27727, 28126, 31015, 30159, 31635, 30958, 29537, 28185, 25355, 23044, 
    21355, 16214, 13031, 7238, 4283, 188, -4482, -8835, -12710, -16777, 
    -20002, -24849, -24727, -26487, -30735, -31393, -31185, -29607, -29905, 
    -26896, -26474, -22363, -19637, -16790, -13591, -10078, -5878, -547, 
    4081, 7007, 12949, 16424, 19691, 22906, 26365, 26493, 29457, 30375, 
    30776, 30805, 28915, 28572, 26172, 24019, 19669, 17840, 13481, 8789, 
    5052, 811, -3736, -8701, -11769, -15925, -18874, -22526, -25019, -28961, 
    -28624, -31522, -29957, -30142, -29964, -28533, -26678, -23923, -20902, 
    -16610, -13853, -9318, -4662, -1397, 2471, 7516, 12401, 14900, 19872, 
    22366, 25039, 28023, 29059, 30153, 31030, 29522, 30053, 27272, 26447, 
    23107, 20038, 18537, 13226, 8536, 6986, 1306, -2495, -8738, -11145, 
    -14857, -19203, -22783, -25647, -26490, -28346, -31233, -31896, -29757, 
    -28368, -29866, -24899, -25689, -21070, -16686, -13950, -9437, -5639, 
    -1354, 2074, 7880, 12261, 14944, 18949, 22351, 25183, 28630, 28796, 
    31051, 32137, 30147, 28948, 29055, 28548, 24704, 21975, 18829, 14313, 
    10856, 4571, 696, -1510, -7419, -11945, -14761, -18748, -21539, -25065, 
    -28410, -30075, -29637, -32116, -30068, -30657, -26803, -27281, -24643, 
    -21867, -18404, -13857, -11212, -6753, -1843, 1492, 7254, 11022, 15160, 
    18690, 22265, 24593, 27503, 28933, 29637, 30676, 31555, 29896, 28942, 
    27791, 25032, 20414, 19796, 13171, 9385, 7382, 615, -2313, -7305, -10169, 
    -14590, -19481, -22322, -25131, -27143, -28473, -31649, -30362, -30734, 
    -29591, -27513, -26893, -25419, -22934, -19014, -14339, -11784, -7294, 
    -1761, 1691, 7554, 11652, 14593, 18098, 20978, 25054, 27543, 29148, 
    29829, 30107, 31354, 30529, 28927, 26833, 25212, 22308, 18910, 15504, 
    10298, 6625, 3563, -1546, -6811, -10234, -14266, -17513, -21744, -24722, 
    -28121, -27439, -29087, -31923, -31686, -29124, -29146, -27459, -24553, 
    -22005, -18979, -14931, -9815, -7566, -2381, 2675, 6863, 10739, 14158, 
    18362, 22373, 23884, 25607, 30064, 29483, 30871, 30188, 29645, 28934, 
    26282, 26355, 21915, 18975, 15715, 10391, 7278, 2908, -1331, -6089, 
    -11798, -14483, -18839, -20723, -25496, -25775, -28130, -30840, -31513, 
    -30010, -29986, -30029, -26753, -26332, -21387, -20077, -16278, -11114, 
    -7120, -3020, 1604, 3985, 10473, 13665, 17568, 20965, 24485, 27513, 
    28464, 29834, 31698, 31699, 30699, 28977, 26469, 24178, 22266, 19093, 
    14719, 11618, 7284, 3475, -702, -5617, -8681, -15056, -18590, -22580, 
    -22569, -26673, -29116, -29392, -30681, -30933, -31323, -28732, -27716, 
    -24114, -21323, -18154, -15215, -11442, -9289, -3037, 2120, 6436, 8756, 
    14208, 18572, 20083, 24980, 25656, 29526, 28880, 30403, 30346, 31180, 
    30789, 28737, 24507, 21137, 18740, 17837, 11813, 7339, 2804, -1108, 
    -5273, -9713, -11806, -17737, -19965, -22912, -26478, -28994, -30017, 
    -30470, -30127, -30853, -29475, -28648, -26874, -23562, -19688, -15858, 
    -12825, -8724, -4298, -168, 4873, 8279, 12297, 16905, 20393, 21944, 
    24707, 27445, 29846, 30037, 29808, 30952, 29294, 26532, 25243, 23772, 
    19435, 16636, 12420, 8539, 4954, -746, -5837, -9484, -13367, -16932, 
    -19206, -23409, -26275, -27507, -29933, -32284, -31496, -29410, -28554, 
    -27514, -24005, -21810, -19975, -15922, -13154, -8566, -4424, 382, 3421, 
    7592, 12912, 17385, 19621, 23354, 26013, 28364, 29715, 30945, 31768, 
    30386, 28828, 29049, 27028, 23993, 20070, 16960, 12120, 9535, 4659, 
    -1059, -5150, -8199, -13773, -16678, -20423, -24386, -26048, -29130, 
    -29038, -29571, -30455, -30136, -30417, -28656, -26438, -23754, -20665, 
    -16861, -13780, -10892, -6073, 73, 2875, 7264, 11014, 17190, 19545, 
    22179, 25145, 28086, 28661, 30116, 31984, 29949, 29744, 28013, 25881, 
    23729, 21480, 17865, 13605, 9056, 4050, -79, -4471, -8683, -12197, 
    -16035, -19522, -24191, -24495, -27682, -29462, -31064, -30732, -32336, 
    -29266, -28646, -24640, -23059, -20575, -16968, -13936, -9600, -5314, 
    -931, 2819, 7774, 11411, 15629, 18912, 21972, 26399, 26252, 29278, 29756, 
    31413, 31252, 30045, 28130, 26786, 24816, 20814, 19221, 12345, 9846, 
    5564, 2043, -3673, -8052, -11775, -15710, -18441, -22030, -25136, -26404, 
    -29796, -30093, -30579, -29700, -29976, -27859, -26822, -24310, -20585, 
    -16666, -13496, -10983, -3825, -1438, 1362, 6907, 11218, 15705, 19456, 
    21148, 25769, 28346, 29482, 29842, 31311, 31783, 30460, 28459, 25645, 
    24227, 20959, 17177, 14039, 8560, 4365, 931, -2742, -7345, -11138, 
    -13847, -20342, -23242, -25435, -27458, -29498, -28802, -30823, -32333, 
    -30656, -28946, -25681, -23737, -21280, -18420, -14206, -10082, -6028, 
    -2559, 2120, 6400, 10995, 15424, 17849, 22058, 24490, 27805, 28535, 
    29888, 31728, 30805, 31235, 28551, 27719, 26285, 21996, 18568, 14643, 
    10404, 5549, 940, -1814, -6105, -12006, -15903, -17506, -21722, -25829, 
    -25759, -27973, -29823, -29818, -29023, -30963, -29943, -27860, -25430, 
    -22958, -17432, -15604, -12235, -6976, -1806, 3243, 6413, 11778, 14191, 
    18516, 22067, 24634, 26498, 28717, 30244, 31467, 28964, 28436, 30240, 
    26667, 25255, 21887, 19859, 14911, 10265, 7821, 2347, -1728, -5226, 
    -11688, -13939, -16641, -21718, -23702, -26644, -28017, -30359, -30532, 
    -31627, -31153, -27617, -27499, -24972, -22306, -20028, -15325, -10408, 
    -7958, -1269, 1510, 7325, 9697, 14840, 18782, 21649, 24186, 27517, 28706, 
    30955, 29481, 31256, 31168, 29199, 27841, 24359, 22485, 20576, 14994, 
    12217, 8067, 1684, -1131, -6387, -9702, -14953, -18043, -21231, -23392, 
    -25134, -28091, -30365, -30633, -30534, -29727, -29029, -26933, -24681, 
    -21178, -19774, -15686, -11598, -7309, -2679, -209, 5180, 9525, 13495, 
    16833, 22277, 25281, 25525, 28156, 30133, 29711, 32067, 31629, 29367, 
    28307, 25178, 23441, 20714, 16346, 11629, 7377, 3225, -1884, -4197, 
    -10961, -13361, -16608, -21175, -23356, -26531, -28678, -29570, -30545, 
    -30300, -31224, -28636, -28731, -25990, -22266, -18782, -15238, -13198, 
    -9201, -4913, 468, 6110, 10552, 14225, 17274, 19946, 22481, 25797, 29831, 
    29620, 29838, 30772, 29128, 29652, 27495, 24315, 23353, 19599, 17299, 
    11750, 6875, 4721, 612, -6047, -10040, -14485, -16939, -19464, -25213, 
    -26637, -27484, -28852, -30352, -31353, -31222, -28624, -28198, -26225, 
    -23324, -20338, -16348, -10928, -7650, -3915, 271, 3310, 7503, 12122, 
    16728, 21516, 21683, 25817, 29605, 30458, 30979, 31344, 30275, 29596, 
    27637, 27070, 24343, 20094, 17882, 12626, 8888, 4045, 1342, -5795, -8953, 
    -13821, -15902, -21144, -23817, -25544, -28689, -30154, -29093, -31623, 
    -30951, -30560, -27764, -27509, -23517, -20090, -15753, -13097, -7947, 
    -4751, 202, 6050, 8479, 12794, 16200, 21712, 23561, 25568, 27347, 29791, 
    29365, 29785, 31213, 30666, 27895, 25674, 24482, 20653, 16368, 13097, 
    7904, 3397, 198, -2635, -8211, -11789, -14816, -19856, -23108, -26336, 
    -27471, -29141, -30414, -30584, -31024, -29491, -28512, -24788, -22508, 
    -21030, -17019, -14540, -9696, -5046, -594, 4019, 7691, 12544, 17383, 
    20451, 22046, 25660, 27602, 28973, 30880, 30247, 30431, 29291, 27710, 
    25580, 23327, 22446, 18956, 14289, 10216, 5246, 498, -2973, -8075, 
    -13411, -16591, -18646, -23267, -24572, -28017, -29675, -31186, -29923, 
    -31485, -29906, -28052, -25429, -23895, -19808, -18168, -13774, -9772, 
    -6044, -1708, 5060, 8260, 11057, 16525, 18302, 21792, 24978, 26192, 
    29509, 30117, 31489, 29460, 30774, 27730, 26598, 23099, 20449, 15904, 
    14833, 10301, 3906, 1131, -3335, -6427, -12937, -15558, -20177, -21988, 
    -25445, -27044, -29667, -30051, -30772, -30396, -29139, -28581, -26553, 
    -23601, -20754, -19286, -15129, -11604, -4794, -786, 2465, 5645, 11975, 
    15334, 17284, 22084, 25612, 27406, 30450, 29777, 30370, 31127, 29700, 
    28317, 26858, 25470, 21245, 17452, 13361, 9488, 5774, 1888, -2935, -8768, 
    -11973, -15017, -19358, -22051, -24538, -26975, -28767, -30637, -31466, 
    -30677, -30407, -27931, -27835, -25954, -23175, -18900, -13833, -9664, 
    -6196, -3045, 3934, 7530, 11310, 15820, 19257, 21652, 23709, 27687, 
    29210, 30408, 30654, 31477, 28712, 27535, 26290, 23993, 21489, 19267, 
    14415, 10807, 6329, 484, -3102, -7611, -10923, -14158, -19805, -21888, 
    -25942, -26258, -28775, -29685, -29636, -31909, -29132, -28613, -27297, 
    -23317, -22714, -18646, -14660, -11387, -6416, -2134, 1790, 6552, 12574, 
    14669, 19901, 21060, 25097, 26028, 29651, 29395, 31927, 30686, 31543, 
    28422, 27666, 25189, 22802, 17958, 14436, 11416, 7453, 2720, -1383, 
    -5132, -10595, -14908, -17704, -22195, -23977, -25734, -28709, -30956, 
    -30651, -30363, -30848, -27897, -27303, -24811, -21018, -18711, -14107, 
    -10970, -7869, -2289, 990, 6991, 10344, 14607, 17801, 22654, 25426, 
    26121, 28316, 31121, 31610, 31774, 31677, 28228, 27445, 24445, 22845, 
    18302, 16418, 12020, 7061, 3009, -1660, -7128, -10440, -13724, -17314, 
    -21358, -24250, -25761, -28127, -28500, -31254, -31201, -30708, -29763, 
    -27445, -25263, -22242, -19558, -16113, -12257, -7489, -4030, -2, 6256, 
    10258, 13912, 17190, 20319, 24840, 26341, 29322, 31363, 30370, 31104, 
    31617, 28591, 27518, 24203, 21488, 20586, 14913, 12227, 7687, 3266, 482, 
    -5824, -9189, -13285, -17741, -21086, -24378, -27722, -28997, -29309, 
    -30907, -31993, -30419, -30125, -27618, -25164, -22300, -20292, -17161, 
    -11303, -6848, -3976, 2288, 5050, 9652, 12932, 16600, 21787, 22693, 
    24805, 29616, 28430, 29296, 29743, 30563, 29656, 27012, 24425, 22570, 
    21028, 17493, 13154, 9021, 4131, -1089, -5908, -9900, -13329, -17750, 
    -20868, -24370, -26293, -28335, -29786, -31964, -32009, -30396, -29758, 
    -27704, -25864, -23830, -19414, -15204, -12429, -9163, -2915, 148, 5367, 
    8812, 14282, 16475, 19906, 23462, 25893, 27069, 29921, 30451, 30751, 
    31054, 29539, 27229, 26200, 21598, 19521, 17127, 11817, 7744, 5396, 320, 
    -4415, -7950, -13588, -17124, -18754, -23867, -25530, -26862, -29645, 
    -30597, -30310, -30169, -30211, -27746, -27185, -22539, -19990, -17102, 
    -13717, -9028, -2662, 738, 4148, 8137, 12824, 16572, 19827, 22737, 26826, 
    28084, 29829, 31126, 32087, 29574, 29143, 28332, 25140, 22086, 19093, 
    16551, 14425, 10476, 5972, -1437, -4133, -8725, -13367, -16601, -20381, 
    -21831, -26268, -28461, -28797, -29603, -30162, -31213, -28254, -28584, 
    -27471, -23138, -19715, -17421, -12392, -9821, -3473, -798, 3913, 8696, 
    12404, 14831, 19024, 21856, 25167, 27503, 29893, 29242, 30695, 29976, 
    28718, 27457, 27605, 24228, 19058, 17177, 12295, 9328, 5294, -967, -4172, 
    -6866, -11578, -16338, -19346, -22546, -25699, -26490, -28603, -30310, 
    -30358, -30573, -30278, -29121, -27995, -24702, -20934, -18517, -14571, 
    -8565, -5753, -111, 3478, 8425, 12917, 17393, 17939, 22664, 25814, 26916, 
    29341, 30257, 29984, 31183, 29743, 29979, 27585, 24716, 19349, 17211, 
    13632, 9410, 6193, -231, -2684, -6863, -11166, -14859, -20811, -22652, 
    -25170, -27499, -27805, -30793, -30579, -30495, -30219, -29892, -26217, 
    -23995, -21691, -18072, -14443, -8494, -6480, -1803, 3761, 7540, 10514, 
    15133, 20426, 21726, 26132, 27187, 29701, 30211, 31294, 29927, 30527, 
    29180, 25838, 23876, 20468, 17086, 14572, 9251, 5611, 1261, -2018, -7178, 
    -10405, -16275, -18961, -22019, -24904, -28827, -30571, -30426, -31457, 
    -31060, -30738, -29331, -26994, -25109, -20884, -16556, -14690, -10707, 
    -5807, -3064, 3341, 7647, 12852, 14079, 18159, 23550, 23931, 28302, 
    29408, 31359, 30670, 30781, 29066, 30123, 25239, 24516, 22962, 16612, 
    14438, 9842, 6232, 2157, -2672, -6245, -12176, -14652, -19643, -21471, 
    -25005, -27742, -27848, -31013, -31221, -31087, -29915, -28326, -27081, 
    -24327, -21941, -17376, -16356, -10209, -6370, -3073, 1338, 6463, 11115, 
    14863, 17296, 22184, 24946, 26766, 29601, 30104, 30744, 32406, 31255, 
    30308, 27567, 24481, 22506, 17495, 14969, 11575, 8164, 2242, -1660, 
    -7008, -10402, -15801, -16840, -21012, -25024, -27205, -27766, -30640, 
    -30589, -31455, -31732, -29397, -27329, -24617, -23405, -19772, -14993, 
    -11872, -7271, -3179, 1748, 5681, 9852, 14967, 18050, 21215, 24573, 
    26127, 29690, 31646, 30711, 30761, 29476, 28961, 25939, 24252, 22013, 
    19508, 15176, 10653, 7924, 3014, -2991, -6405, -10034, -12914, -18232, 
    -22431, -23999, -26554, -28241, -29673, -30400, -31139, -29844, -28629, 
    -25911, -25369, -21646, -18005, -16741, -11886, -8243, -3641, 1718, 6660, 
    9685, 14393, 17048, 22185, 24103, 25637, 28297, 29160, 31398, 29649, 
    29271, 30042, 27831, 24354, 23815, 20103, 15418, 12548, 8599, 3862, 
    -1438, -6702, -10545, -15149, -16811, -20716, -24878, -26293, -28907, 
    -29467, -31641, -31503, -28759, -29411, -27623, -24241, -21842, -20476, 
    -16021, -10821, -8495, -2844, 751, 5650, 8951, 13058, 17023, 20300, 
    23145, 25909, 27569, 29146, 30101, 29351, 30824, 29196, 29046, 24219, 
    21355, 19322, 15181, 11898, 8138, 3601, 157, -4003, -9413, -14518, 
    -17418, -19279, -23874, -25582, -28029, -29617, -30168, -31379, -30530, 
    -29514, -28362, -25361, -22223, -18793, -16485, -11581, -7950, -2812, 
    1617, 6013, 8773, 13561, 18498, 21013, 23215, 26323, 27310, 29638, 30522, 
    30369, 31355, 29375, 27999, 26382, 21492, 20375, 16175, 12756, 8539, 
    3472, -1612, -4453, -7963, -11562, -17097, -20415, -23628, -26055, 
    -27623, -29586, -29365, -32319, -29690, -29988, -27336, -24665, -22147, 
    -19521, -17436, -12062, -9017, -5465, 1087, 2746, 7905, 13702, 16822, 
    19219, 25034, 25831, 28339, 29019, 30799, 30816, 30904, 30710, 27864, 
    26616, 21619, 21942, 17204, 13356, 8995, 3801, 2089, -3998, -8038, 
    -12351, -15110, -20121, -23535, -26393, -27453, -30815, -30003, -30757, 
    -30059, -30952, -28056, -24890, -24809, -22005, -18275, -13820, -9085, 
    -5528, -401, 5404, 8762, 12173, 16229, 18761, 23365, 25224, 27575, 30479, 
    28570, 31107, 29852, 29622, 28500, 26857, 23222, 21637, 18240, 13716, 
    8292, 4092, 1953, -3605, -7169, -12393, -15653, -18951, -22226, -25166, 
    -27243, -29594, -30274, -30078, -30951, -29831, -28205, -25768, -24902, 
    -21928, -17547, -13710, -9084, -5245, 719, 4146, 7412, 11765, 16170, 
    20358, 22772, 25016, 28211, 28486, 31380, 32338, 29849, 31033, 27627, 
    26322, 23572, 20957, 16250, 15003, 8630, 4552, 1796, -3610, -7866, 
    -12088, -15506, -19752, -22470, -26097, -27459, -29875, -30213, -31790, 
    -29399, -29780, -29388, -26399, -25910, -19260, -18343, -15516, -10853, 
    -6313, -1511, 3365, 6413, 12423, 14689, 18764, 23716, 26730, 27989, 
    29744, 31604, 30290, 32313, 30966, 27346, 25681, 24438, 20005, 18028, 
    14483, 9282, 5192, 792, -2424, -7927, -11316, -15510, -18113, -21009, 
    -24393, -26691, -29332, -28830, -31076, -30650, -31094, -27942, -26126, 
    -24842, -20853, -16695, -14765, -9165, -6145, -790, 2294, 7712, 11548, 
    15156, 18892, 21791, 23998, 26454, 28987, 31424, 30323, 30604, 29723, 
    28493, 26920, 24732, 21458, 19493, 15572, 11391, 6392, 2414, -1555, 
    -6815, -10334, -15008, -18577, -22217, -24634, -27271, -29268, -31443, 
    -32280, -29988, -30902, -29572, -27880, -24676, -22138, -17632, -15204, 
    -11461, -8244, -1891, 2400, 7017, 11610, 15068, 18371, 22002, 24253, 
    25882, 28969, 30401, 30691, 30884, 29060, 28415, 26838, 24372, 20429, 
    19503, 16008, 10648, 7041, 3453, -3354, -6680, -11147, -14580, -18273, 
    -21131, -24184, -25852, -27468, -30288, -29862, -31973, -31102, -29458, 
    -26423, -25901, -22362, -18731, -14622, -9459, -5850, -1787, 2587, 7115, 
    9780, 15707, 18830, 21474, 23288, 27825, 28882, 30041, 30628, 29703, 
    30793, 29909, 27581, 25675, 23024, 19552, 14966, 10843, 8001, 3941, 
    -1450, -6070, -11625, -13401, -18268, -21971, -24290, -27786, -29079, 
    -28368, -30690, -31295, -31239, -29807, -28210, -24373, -22812, -19369, 
    -14490, -11522, -6890, -4248, 1699, 5435, 10396, 13841, 17195, 22772, 
    24047, 25300, 29778, 30101, 30189, 31949, 31056, 30251, 27237, 24580, 
    21623, 19124, 13867, 11676, 9274, 2969, -856, -5819, -9767, -12936, 
    -17899, -22147, -24172, -27009, -26837, -30764, -30137, -31036, -29648, 
    -28712, -27008, -27145, -23575, -20796, -16486, -13304, -8880, -3870, 
    548, 4448, 9723, 14308, 16001, 21465, 23829, 27512, 29780, 30251, 31534, 
    31352, 31541, 29160, 29387, 24687, 22171, 20247, 14755, 11623, 8619, 
    3737, -1600, -5690, -8513, -13351, -17372, -20068, -25326, -27211, 
    -28460, -28635, -31463, -30333, -30906, -30899, -28607, -26048, -22736, 
    -20808, -15624, -11631, -7347, -3613, 1503, 6031, 9404, 12974, 17610, 
    20407, 22367, 25812, 28536, 29301, 30019, 31343, 30833, 30458, 26903, 
    25548, 22386, 19928, 16232, 12278, 7468, 4535, -363, -3450, -9338, 
    -12328, -16953, -21521, -22693, -24650, -28128, -30364, -30656, -31949, 
    -30453, -29786, -29368, -26145, -23833, -20619, -15221, -13077, -8627, 
    -3646, 1754, 5355, 8029, 14157, 16040, 20224, 21677, 25215, 29235, 29757, 
    30065, 30429, 30804, 29628, 28029, 26030, 24476, 19584, 16709, 12446, 
    8552, 4760, 1587, -4141, -8288, -14113, -14712, -21246, -23543, -26402, 
    -27079, -29056, -30947, -30901, -30789, -30848, -28276, -26115, -22421, 
    -20515, -17131, -11872, -8176, -4348, -287, 3715, 7764, 12632, 15508, 
    19019, 23448, 26887, 26542, 28320, 31382, 30398, 30853, 30058, 27530, 
    25235, 24030, 20366, 17139, 13480, 9199, 4630, 1640, -4584, -8054, 
    -11813, -16404, -19983, -22128, -24422, -27447, -28808, -30578, -30784, 
    -30955, -28837, -27859, -26292, -24219, -19914, -18238, -13043, -10169, 
    -5828, -1027, 3368, 6904, 12027, 15431, 19383, 22080, 25642, 27076, 
    29192, 30261, 30458, 29444, 29617, 27913, 26830, 23702, 19971, 17459, 
    14347, 9644, 6354, 509, -3624, -9158, -12966, -14742, -20635, -23409, 
    -24490, -26596, -28732, -30504, -31428, -30106, -30172, -29726, -27522, 
    -24855, -21772, -17208, -15216, -8716, -6058, -1814, 3864, 7479, 11667, 
    14405, 19345, 22493, 26438, 28593, 27752, 32040, 30581, 30987, 30098, 
    27119, 25391, 25032, 20603, 16423, 14031, 11186, 7043, 625, -3151, -7433, 
    -11152, -15807, -19080, -22588, -25134, -27500, -28826, -28976, -32583, 
    -31551, -31116, -28660, -26575, -23176, -20007, -17799, -13315, -10377, 
    -5271, -2060, 1747, 6820, 12366, 15604, 20360, 22471, 25376, 27836, 
    28735, 30043, 32433, 30840, 30610, 29033, 27262, 23655, 20921, 18708, 
    13414, 11875, 4728, 2082, -1825, -7558, -10577, -15395, -18798, -22021, 
    -24225, -26269, -28562, -30203, -30320, -31761, -29493, -28584, -27613, 
    -23336, -22372, -19074, -13443, -10525, -5044, -2577, 1435, 6146, 10047, 
    14245, 19229, 21719, 25198, 25952, 28933, 30684, 30103, 30949, 30192, 
    28261, 26204, 23474, 23023, 18252, 14759, 11453, 7807, 1973, -2903, 
    -5982, -10325, -14751, -18760, -21431, -24127, -27388, -27901, -30189, 
    -29477, -31216, -29095, -27902, -26934, -23806, -23295, -19692, -15190, 
    -11005, -7857, -3544, 378, 6991, 10294, 13689, 17061, 22678, 25042, 
    27612, 28577, 29485, 31425, 29706, 29978, 29399, 27164, 25068, 21483, 
    19924, 16805, 11912, 7043, 2987, -1153, -5419, -10493, -13427, -17377, 
    -20271, -23726, -26377, -28812, -30267, -31305, -30197, -29047, -28657, 
    -27345, -26271, -21905, -18812, -15802, -11068, -7420, -4921, 883, 5207, 
    9342, 13850, 17996, 21113, 23312, 26008, 28612, 29377, 30242, 30781, 
    30946, 28885, 26796, 25288, 22979, 18008, 17132, 11744, 7354, 3990, 
    -1373, -4566, -9054, -12378, -16892, -20547, -22601, -27950, -29454, 
    -29724, -31323, -30904, -29189, -28680, -27767, -25604, -23042, -19413, 
    -16790, -12397, -8642, -3460, 2085, 3920, 9585, 12739, 15808, 21514, 
    23948, 26251, 27489, 29353, 30659, 30071, 31204, 29412, 28465, 26079, 
    22677, 20787, 16033, 11360, 8577, 3759, -457, -5806, -8964, -13641, 
    -18595, -20434, -23752, -25767, -28635, -30595, -31285, -32274, -30133, 
    -27833, -28867, -25578, -23221, -20444, -15480, -12954, -7260, -3808, 
    1094, 4612, 9325, 13338, 16937, 20872, 24716, 27482, 27201, 30140, 31927, 
    31334, 30560, 28586, 27643, 25318, 22899, 20269, 15952, 12194, 7112, 
    4211, 894, -5902, -8241, -14672, -16533, -20036, -23190, -27389, -28737, 
    -29319, -30215, -31121, -29896, -30849, -27515, -25912, -24272, -21124, 
    -16455, -12985, -8846, -2869, -481, 5494, 7588, 14436, 16384, 21164, 
    24459, 25853, 29106, 29644, 30350, 30220, 30730, 30412, 27887, 26617, 
    24084, 19717, 18548, 11427, 8764, 3430, -402, -4661, -8035, -10931, 
    -17000, -19840, -23345, -25280, -27524, -28331, -31512, -31537, -30756, 
    -31212, -27271, -27307, -24164, -21835, -16332, -11782, -9414, -3840, 
    -231, 3296, 8448, 12665, 15907, 19939, 24013, 24810, 27321, 29602, 30403, 
    30875, 31144, 31050, 29132, 27239, 24984, 21806, 17342, 13740, 9986, 
    3775, 823, -2427, -9504, -12585, -15742, -19677, -23646, -26623, -27901, 
    -30633, -29151, -29502, -29087, -30531, -27990, -27220, -23849, -21617, 
    -18095, -14644, -9552, -5424, -1056, 2314, 7384, 11792, 16412, 19881, 
    22770, 25450, 26897, 28125, 30126, 30948, 30133, 31266, 29104, 26934, 
    24330, 22152, 17122, 15342, 9734, 5861, 938, -3901, -7310, -11150, 
    -16470, -18163, -23225, -25299, -28719, -30980, -31275, -31042, -29017, 
    -29224, -27572, -25886, -22926, -21978, -18792, -15089, -9610, -5164, 
    -280, 3565, 8232, 12114, 15756, 18429, 20567, 24171, 28466, 29232, 29322, 
    29449, 31432, 30934, 28138, 26544, 23933, 21771, 17853, 14743, 9190, 
    5978, 3019, -3004, -8848, -10728, -14866, -20381, -22189, -26843, -27744, 
    -28920, -29898, -30032, -29344, -31302, -30014, -26949, -25534, -21481, 
    -19031, -14430, -11209, -7151, -634, 3158, 8565, 11022, 15721, 20254, 
    21051, 25371, 27953, 28609, 31465, 32161, 30770, 28863, 29613, 26151, 
    25479, 21577, 17548, 15249, 10967, 6607, 2710, -1249, -7334, -11205, 
    -14181, -18879, -21415, -25278, -27048, -28719, -29354, -31209, -30400, 
    -30200, -30643, -26954, -23377, -20516, -17442, -14669, -9502, -4926, 
    -2277, 1848, 7910, 10841, 12985, 18127, 20935, 24536, 27467, 29958, 
    29559, 29374, 31146, 29910, 28252, 26589, 24910, 20258, 18551, 15337, 
    12046, 7025, 2752, -1363, -5892, -9359, -16048, -17872, -22842, -23211, 
    -27219, -28100, -30558, -30898, -29708, -30090, -29037, -28629, -25902, 
    -22685, -17291, -15747, -11206, -7648, -3098, 2438, 7698, 8711, 14886, 
    18035, 22102, 23845, 26266, 29764, 30395, 31422, 30373, 30253, 29007, 
    26630, 25721, 23351, 19693, 16003, 9777, 7022, 3714, -1374, -5228, 
    -10227, -15667, -17130, -20528, -25194, -25947, -28881, -31302, -31281, 
    -29807, -30730, -28826, -27444, -24873, -23075, -18012, -17165, -10349, 
    -6500, -3361, 860, 6851, 9294, 13837, 17131, 19904, 23994, 26777, 28792, 
    29711, 31840, 31495, 29360, 28580, 27412, 24601, 22664, 19677, 15989, 
    11327, 8189, 3940, -857, -5350, -9756, -14970, -17747, -19403, -23802, 
    -24887, -28610, -30905, -31795, -31013, -30305, -30207, -27816, -25514, 
    -22255, -20845, -16209, -13104, -7641, -3084, 111, 6597, 9786, 13785, 
    16221, 20119, 23308, 26543, 27545, 29651, 30266, 31314, 31766, 29442, 
    28635, 25701, 23804, 19921, 16229, 11516, 6958, 2904, -1822, -3926, 
    -9085, -12952, -16709, -21461, -23121, -27250, -28283, -29538, -30784, 
    -30489, -30707, -28775, -28698, -25658, -23300, -19406, -16382, -10608, 
    -7358, -3796, 359, 3123, 9711, 13399, 18119, 20437, 24117, 27165, 29021, 
    28514, 31555, 31765, 30875, 30086, 28153, 25299, 22687, 21129, 16035, 
    12946, 8517, 4086, -388, -4847, -9831, -13975, -15568, -20225, -23852, 
    -24270, -26911, -29964, -31473, -29579, -29677, -30392, -29091, -26483, 
    -23447, -19900, -16871, -12548, -10447, -2973, 235, 5038, 10511, 12077, 
    15831, 18679, 23128, 25256, 27354, 29444, 30790, 31372, 29201, 28367, 
    26918, 27055, 22384, 21297, 16577, 12579, 9151, 3742, -306, -3911, -9903, 
    -11287, -15988, -19008, -22509, -24870, -28259, -30059, -30980, -31913, 
    -30928, -29596, -28210, -26252, -23738, -20998, -16131, -13194, -8278, 
    -4557, -419, 5624, 6878, 11639, 17170, 18584, 22669, 26266, 27093, 29221, 
    30845, 29809, 30909, 28279, 27569, 25683, 22250, 19066, 16103, 13122, 
    9203, 4478, 247, -2248, -7536, -13800, -15792, -18575, -22760, -25592, 
    -28615, -29411, -31158, -32274, -31448, -29343, -28082, -26168, -23604, 
    -21410, -15915, -14270, -9818, -4642, -2172, 3185, 6747, 11625, 16393, 
    19555, 22024, 24730, 27008, 29876, 30322, 31993, 29987, 30659, 28709, 
    27077, 24090, 20478, 16322, 14474, 9977, 6928, 1918, -2719, -7793, 
    -13096, -15193, -20821, -23935, -25696, -28371, -28640, -28558, -31220, 
    -30643, -30118, -28856, -25096, -23697, -20186, -18066, -13355, -10933, 
    -4898, -340, 1523, 6110, 10007, 15914, 19532, 23820, 24895, 26708, 28434, 
    30420, 30299, 30977, 29269, 28369, 27121, 24206, 19987, 18609, 14412, 
    10191, 4856, 2813, -2912, -6202, -11156, -15756, -19355, -21673, -25275, 
    -26616, -29196, -30160, -30754, -30268, -29231, -28476, -26397, -23391, 
    -21370, -17867, -14112, -10846, -7026, -1191, 2074, 6100, 11154, 14469, 
    19321, 22443, 23903, 26975, 29503, 29673, 31000, 30332, 29685, 28935, 
    26962, 24409, 19845, 17744, 14611, 11611, 5037, 2451, -2242, -5928, 
    -11675, -13990, -19704, -22675, -23838, -25906, -29772, -30688, -30497, 
    -30956, -28423, -28692, -25829, -24585, -21645, -19268, -13720, -9622, 
    -5749, -1699, 3409, 6254, 9982, 14240, 18654, 23073, 23650, 25695, 30175, 
    29855, 31619, 32307, 30799, 28010, 28332, 25055, 21798, 18526, 14535, 
    10658, 7770, 1363, -1741, -6283, -9891, -14896, -19190, -21045, -23257, 
    -25878, -29004, -29299, -30140, -29213, -30249, -29867, -27152, -26296, 
    -21820, -19521, -16029, -10038, -7580, -2842, 208, 7029, 10630, 15829, 
    17612, 21332, 24663, 26942, 29690, 31683, 30857, 31273, 29148, 28188, 
    28417, 25351, 22174, 18827, 16490, 10839, 6347, 2133, -2408, -5325, 
    -10137, -14868, -18404, -21804, -23464, -25113, -28696, -31212, -30484, 
    -30471, -31081, -28241, -27089, -23599, -21270, -19528, -16052, -10219, 
    -7285, -3920, 1180, 4044, 9652, 14678, 17538, 21359, 25335, 28161, 28906, 
    30031, 30235, 30515, 30520, 28890, 27818, 25146, 22054, 19404, 14641, 
    11440, 7413, 2191, -161, -4874, -10802, -14263, -17597, -20147, -24421, 
    -27385, -27770, -30387, -31033, -29571, -30145, -29210, -28027, -26502, 
    -22603, -21115, -16059, -12316, -7626, -3225, 1824, 5162, 9804, 12586, 
    17607, 22272, 24543, 26325, 29280, 30040, 31382, 31372, 29993, 29333, 
    28318, 26213, 21390, 19583, 16594, 13158, 8093, 3597, -687, -4373, -9261, 
    -14891, -17459, -20073, -24719, -26997, -28406, -29604, -30066, -30612, 
    -31266, -28062, -27846, -24893, -21257, -20861, -14920, -12206, -8452, 
    -5002, -555, 4322, 8110, 13154, 18648, 19697, 23789, 25545, 27485, 29715, 
    30888, 31613, 30352, 29116, 28228, 27222, 24295, 20266, 15896, 11641, 
    7597, 4869, 172, -4936, -7245, -12160, -16494, -20476, -22584, -25727, 
    -29022, -29945, -30979, -30355, -31495, -30065, -27746, -25873, -22800, 
    -21946, -15443, -13044, -7978, -3580, -104, 3493, 8684, 12865, 16796, 
    20432, 23037, 26684, 27014, 29212, 30219, 31103, 28927, 28271, 26956, 
    26010, 22497, 20596, 16526, 13824, 8636, 3963, 604, -4171, -7016, -12983, 
    -16652, -19184, -23221, -26900, -27497, -28534, -31639, -29324, -31607, 
    -30216, -28882, -27443, -21834, -21187, -18595, -14000, -8406, -4930, 
    536, 4965, 7868, 13088, 16084, 19674, 23808, 26248, 27942, 29952, 31542, 
    31139, 31148, 30766, 29085, 27181, 24912, 19979, 18031, 12993, 8634, 
    4677, -185, -5095, -7988, -11409, -15839, -19445, -23311, -26100, -26789, 
    -30356, -29800, -29777, -29576, -30433, -27560, -27654, -24150, -19897, 
    -16249, -15039, -8451, -3974, -89, 3164, 8034, 12111, 15254, 20539, 
    22104, 26386, 27851, 29361, 29173, 31384, 30581, 29980, 28536, 25913, 
    24570, 21562, 17671, 13881, 9877, 5059, 648, -2207, -5832, -13328, 
    -16473, -19412, -21251, -25658, -27457, -29490, -30888, -30299, -30102, 
    -29992, -28398, -26489, -22720, -21624, -17473, -12482, -9932, -5181, 
    -851, 1260, 7575, 12276, 15512, 18099, 22193, 25036, 26144, 28710, 29700, 
    32115, 31232, 30661, 29194, 26233, 25295, 21617, 17893, 14521, 9766, 
    4764, 2023, -3040, -7559, -11119, -15078, -19597, -22071, -24382, -26493, 
    -29669, -31069, -30572, -31294, -30065, -28821, -26258, -24718, -20660, 
    -18939, -12527, -11269, -6690, -986, 3940, 7911, 11071, 14155, 17926, 
    22738, 24970, 27904, 28812, 30798, 32123, 30493, 29555, 28058, 25827, 
    25130, 21770, 17790, 14828, 9978, 8061, 2523, -3543, -8250, -11282, 
    -13747, -17197, -21434, -25245, -28294, -30362, -29910, -30826, -29330, 
    -30979, -29311, -26672, -24584, -22118, -18564, -16112, -11173, -6305, 
    -1609, 1941, 6390, 11150, 13269, 19154, 21838, 24894, 25862, 29142, 
    30662, 31941, 30769, 30555, 29090, 27491, 24557, 21296, 17683, 14971, 
    11593, 6891, 1567, -2822, -5197, -10061, -14606, -18417, -21234, -24141, 
    -26981, -28882, -29954, -29808, -31387, -29954, -28601, -26220, -24249, 
    -21705, -18001, -13984, -10864, -7982, -3810, 806, 6209, 10464, 14344, 
    18454, 21597, 23642, 26591, 28386, 29171, 30765, 31155, 30195, 29287, 
    26847, 26452, 22542, 19290, 15207, 11616, 8158, 3984, -886, -6695, 
    -10379, -14750, -18235, -20414, -24388, -26109, -26882, -30912, -31029, 
    -30161, -30980, -29051, -25982, -26611, -22887, -19753, -15285, -10974, 
    -7422, -3352, 524, 6407, 11318, 12393, 19331, 20558, 23907, 25680, 28413, 
    30518, 30656, 30319, 29868, 27636, 26740, 25837, 22258, 17692, 15230, 
    10729, 8052, 4659, -748, -4381, -10089, -13338, -17557, -19865, -22551, 
    -27800, -27582, -30220, -30055, -31377, -29925, -28933, -28098, -25625, 
    -23459, -18963, -14442, -10865, -7297, -3356, 1952, 6919, 9512, 12916, 
    17630, 21184, 23811, 25178, 28023, 29804, 30545, 30822, 30081, 29689, 
    27838, 26347, 21878, 19976, 16923, 10805, 8638, 3791, 628, -4387, -8235, 
    -13343, -17575, -21983, -21981, -26206, -27704, -29871, -29490, -29297, 
    -31225, -30728, -26945, -26023, -23953, -19013, -16837, -12300, -9643, 
    -4145, 1046, 3428, 8272, 13394, 15693, 19357, 23531, 25292, 27897, 30239, 
    29468, 31307, 31983, 30265, 28473, 25128, 21759, 20659, 16887, 11953, 
    8719, 4174, -458, -4548, -7868, -14058, -16518, -19066, -23500, -26775, 
    -29274, -30148, -31129, -29355, -30077, -30491, -28005, -26602, -24922, 
    -20392, -16380, -13917, -8738, -3270, 111, 3116, 10307, 13434, 16620, 
    18682, 23690, 25311, 29204, 30706, 29314, 29845, 30635, 30649, 27868, 
    26404, 22724, 21323, 17956, 12948, 7774, 4114, 1408, -3188, -9674, 
    -13815, -16624, -19097, -22414, -25127, -28637, -29673, -30536, -30472, 
    -32022, -31003, -28359, -27308, -22697, -19768, -18282, -13948, -7795, 
    -5793, -862, 4940, 9376, 12800, 16073, 20955, 21288, 25991, 27842, 30331, 
    31252, 30694, 31133, 30052, 28891, 27322, 23210, 20603, 16866, 13136, 
    9457, 5396, 1174, -2568, -7996, -13198, -16055, -19564, -21558, -25354, 
    -27301, -29818, -29605, -31171, -30304, -30162, -26817, -27101, -23194, 
    -21210, -17581, -13407, -10859, -3891, -1705, 4674, 6648, 12800, 14985, 
    20046, 22668, 23682, 27656, 28689, 29743, 31140, 31177, 30170, 28644, 
    26670, 23730, 21189, 18678, 13857, 10965, 7161, 137, -3107, -6802, 
    -12897, -16824, -18665, -21495, -25704, -27723, -29897, -30155, -30351, 
    -30309, -29294, -28693, -26181, -25046, -20681, -17057, -13972, -9380, 
    -5591, -33, 3389, 7133, 11405, 14297, 18621, 22928, 25335, 27849, 29388, 
    29369, 31168, 30388, 29564, 29979, 25302, 24997, 22736, 17649, 15461, 
    9450, 5134, 930, -1964, -6971, -12044, -15746, -17314, -20935, -24234, 
    -27670, -28675, -29987, -30498, -29817, -28330, -29706, -26775, -24647, 
    -20185, -18409, -14364, -10064, -5653, -3322, 3743, 5905, 11455, 16975, 
    19102, 21798, 24172, 27458, 27640, 30095, 30974, 31350, 31137, 29159, 
    26109, 23636, 22062, 18452, 13878, 9848, 5918, 2010, -1830, -5734, 
    -10943, -15283, -19666, -21509, -24915, -28622, -30228, -29106, -29705, 
    -30835, -31203, -27553, -26603, -25543, -22941, -17801, -15019, -10756, 
    -7488, -2609, 1931, 6888, 10887, 15937, 18037, 21528, 23446, 27355, 
    28444, 29533, 31913, 30465, 29695, 28347, 27640, 24877, 22579, 19974, 
    14172, 10883, 5804, 1371, -775, -6311, -10382, -15456, -18581, -21383, 
    -22868, -27207, -28939, -28685, -31680, -32474, -30340, -30101, -28417, 
    -24996, -21289, -19397, -15468, -9836, -8612, -3012, 516, 6169, 9991, 
    14540, 17476, 20397, 24734, 25967, 27334, 30540, 31095, 31616, 30136, 
    30072, 26992, 25638, 21848, 20002, 14463, 11930, 6037, 1732, -58, -6666, 
    -11443, -14006, -18515, -21010, -25059, -26532, -28009, -30496, -30981, 
    -30137, -30521, -29072, -26673, -26300, -22004, -18270, -16068, -12212, 
    -7997, -4221, 1323, 5923, 10388, 13531, 18351, 21300, 25458, 26133, 
    27592, 30860, 31058, 30225, 30143, 29308, 26057, 24318, 21991, 19442, 
    16567, 11649, 8145, 3565, -780, -4290, -9938, -12890, -18065, -21599, 
    -22884, -26649, -29286, -29066, -29805, -30755, -30457, -28631, -27746, 
    -26312, -23495, -20744, -16357, -12490, -8053, -4797, -174, 6470, 9634, 
    15015, 17298, 20408, 23706, 27912, 27811, 29749, 31459, 31783, 29617, 
    30299, 27607, 26213, 22110, 20189, 16727, 13875, 8811, 3461, -1011, 
    -5345, -8875, -13576, -18282, -20171, -23561, -25192, -29438, -29573, 
    -30045, -31578, -30127, -29769, -27868, -26797, -22660, -18559, -17772, 
    -11648, -7383, -3078, 393, 3677, 8954, 12331, 16547, 20593, 22554, 26705, 
    28404, 30246, 31958, 31040, 29902, 29880, 26982, 25124, 21883, 20603, 
    17214, 13616, 7821, 3691, 760, -5170, -9973, -14790, -17852, -20677, 
    -23692, -26296, -28244, -29311, -29659, -30538, -30821, -30704, -28479, 
    -26816, -24168, -19896, -17129, -12842, -9574, -4362, -27, 3370, 8828, 
    12462, 17812, 21072, 22247, 24501, 27922, 29274, 30702, 31507, 30586, 
    29450, 28566, 25315, 22738, 20199, 16093, 13641, 9731, 3771, -247, -4232, 
    -7656, -12672, -16546, -20297, -24129, -24734, -27684, -30735, -31246, 
    -31279, -29839, -29728, -28735, -25336, -24939, -20632, -16154, -13794, 
    -9160, -5325, 429, 4164, 7962, 11357, 15698, 18200, 23555, 27057, 28585, 
    30609, 30112, 31452, 31633, 28984, 28739, 26021, 22702, 21901, 15919, 
    13386, 9496, 5167, 1863, -3179, -8757, -13107, -17212, -19580, -23951, 
    -25513, -27602, -29712, -29683, -31182, -31236, -30466, -28237, -28173, 
    -24416, -20779, -17864, -13275, -9147, -4108, -971, 3113, 7625, 11468, 
    15854, 19404, 22869, 25003, 27753, 30134, 30524, 30767, 29214, 30257, 
    29421, 24939, 24372, 22163, 18339, 12914, 10626, 5766, 1248, -2300, 
    -6103, -11469, -16577, -19448, -22681, -25088, -27686, -27605, -29432, 
    -31234, -31765, -30157, -28280, -26329, -23622, -21987, -17649, -14196, 
    -9898, -5122, -185, 2855, 5771, 11653, 13810, 19680, 22360, 25026, 26357, 
    29747, 31112, 29599, 30487, 29879, 27845, 27036, 24916, 21977, 16286, 
    12508, 9853, 5551, 219, -1435, -6967, -11746, -15999, -18693, -23029, 
    -26122, -28025, -30224, -29270, -30868, -30644, -29758, -27776, -27223, 
    -22780, -21639, -18123, -13549, -10135, -6830, -779, 2673, 6223, 10147, 
    16054, 18450, 22159, 26135, 27173, 29435, 30334, 30355, 30936, 31279, 
    29128, 25693, 25002, 21850, 18695, 13711, 10434, 5948, 1410, -2333, 
    -5672, -11153, -15181, -17790, -20458, -25487, -26212, -29760, -30849, 
    -31035, -32034, -29028, -29368, -28156, -23308, -22965, -19206, -16204, 
    -10396, -7480, -1575, 2716, 5995, 10954, 15946, 18407, 21766, 24598, 
    28695, 30506, 29769, 31476, 32085, 28980, 29228, 28031, 23673, 22114, 
    18410, 14068, 11666, 6735, 3366, -1771, -7199, -10507, -14171, -17355, 
    -20513, -24163, -26643, -29993, -30223, -30001, -30505, -29847, -28556, 
    -27161, -24451, -22345, -18426, -16118, -11135, -7477, -2300, 1892, 5449, 
    10335, 13833, 18067, 20978, 24216, 26311, 28612, 29695, 30418, 31477, 
    29338, 28495, 27304, 24348, 22767, 17876, 14968, 9569, 6370, 3415, -713, 
    -6580, -9543, -13879, -19048, -21588, -23995, -26938, -29201, -29327, 
    -31289, -30035, -30304, -28537, -26562, -24319, -22354, -19448, -14956, 
    -11309, -6384, -1906, 1091, 4365, 9986, 15296, 17431, 20330, 24743, 
    26580, 27683, 30024, 30048, 31626, 31900, 29207, 27257, 24835, 22820, 
    19382, 15410, 12629, 7653, 3931, -2284, -5712, -10456, -13229, -17240, 
    -21554, -23003, -26265, -28818, -28486, -30725, -30442, -30946, -28371, 
    -29274, -25252, -21955, -19749, -15954, -13280, -8196, -3256, 104, 5298, 
    8373, 13380, 17339, 19111, 23421, 26056, 28091, 28793, 30946, 30971, 
    29726, 28715, 27151, 26272, 21098, 18691, 16928, 12356, 9292, 4521, -536, 
    -5378, -10328, -14534, -16420, -19005, -22838, -26345, -27071, -29125, 
    -29241, -31811, -29841, -29087, -27773, -26110, -22754, -18183, -16308, 
    -12660, -7652, -2713, -107, 4779, 9073, 13086, 16370, 20652, 23790, 
    26553, 27943, 29893, 30990, 29917, 30605, 29599, 27658, 26025, 22387, 
    19584, 16385, 11672, 8664, 5374, -752, -5543, -7584, -11877, -16061, 
    -18895, -23123, -25188, -28591, -29212, -30608, -29681, -31730, -28639, 
    -26633, -26682, -22111, -21106, -17539, -13906, -8141, -5485, -1463, 
    3483, 9184, 12598, 15070, 19657, 24605, 26586, 27774, 28932, 30304, 
    30540, 29188, 27966, 28526, 25675, 23673, 20688, 17716, 11973, 7945, 
    4307, 522, -4183, -8980, -11089, -15406, -21166, -24039, -26849, -27351, 
    -28887, -29947, -30144, -30463, -30916, -28584, -24827, -22304, -19823, 
    -16928, -13360, -8993, -4546, 282, 4233, 8627, 13235, 15770, 20126, 
    21844, 24007, 26975, 27770, 31803, 29978, 29174, 28470, 29600, 26830, 
    23194, 21256, 17902, 13341, 10082, 4977, 1975, -4367, -7886, -11328, 
    -16786, -19582, -21645, -24479, -28938, -28794, -29926, -30470, -30784, 
    -30020, -28862, -27677, -24620, -19060, -18838, -13859, -10749, -4723, 
    -1130, 3695, 7323, 11349, 16105, 19772, 21908, 25913, 29467, 29128, 
    29620, 30843, 30021, 29676, 29461, 26475, 23197, 20646, 17742, 12302, 
    10342, 7120, 2934, -4355, -7801, -12410, -15836, -18532, -23100, -24645, 
    -26655, -28934, -30239, -29337, -29804, -29990, -27520, -26435, -23924, 
    -21218, -17404, -14599, -11195, -6470, -771, 3027, 7681, 11183, 15654, 
    19200, 23229, 25043, 27482, 28764, 30072, 29745, 30675, 28406, 29388, 
    27352, 24423, 21183, 18528, 12725, 8794, 6007, 526, -1769, -5490, -10964, 
    -13558, -19226, -23507, -25539, -26727, -29908, -31177, -29809, -30020, 
    -30005, -28618, -27995, -25124, -20836, -18569, -15047, -9660, -5672, 
    -2120, 2479, 8856, 10001, 16256, 18953, 20727, 26206, 27653, 28546, 
    31321, 30617, 30842, 31340, 29047, 26527, 23998, 22774, 18223, 14825, 
    10613, 5053, 1908, -2136, -7685, -10692, -15274, -18053, -20176, -24770, 
    -27329, -28841, -29906, -31112, -29546, -31500, -30198, -26799, -25099, 
    -20902, -19826, -13542, -9856, -7529, -2181, 1357, 6329, 9932, 14065, 
    17994, 21422, 25590, 26050, 29616, 31723, 30337, 29875, 31167, 27553, 
    26735, 24494, 20917, 18848, 15383, 10383, 6522, 1015, -722, -7437, 
    -11713, -14524, -19000, -21534, -23804, -27251, -29382, -30834, -30626, 
    -30285, -30181, -28320, -25793, -24291, -22464, -17691, -14135, -11547, 
    -5965, -4282, 1378, 4622, 11868, 14456, 17565, 22656, 24554, 25520, 
    26980, 29895, 31060, 30956, 30839, 27911, 27853, 25020, 21711, 17786, 
    15213, 10862, 7601, 3421, 183, -5668, -10137, -14357, -19376, -21536, 
    -23134, -27279, -26939, -29258, -30250, -31051, -29920, -29391, -28679, 
    -25176, -22481, -19516, -16437, -10457, -6255, -4132, 1756, 6196, 8851, 
    13383, 18701, 20908, 23529, 27250, 28917, 30139, 30713, 31225, 30396, 
    29318, 27558, 25428, 23363, 20025, 14511, 10196, 7643, 2116, -1256, 
    -5989, -9753, -14143, -17382, -21221, -23794, -26239, -27422, -28549, 
    -31577, -30895, -29928, -29925, -26856, -25377, -23836, -20836, -15660, 
    -12308, -9289, -3618, 1599, 5706, 10079, 13248, 17335, 22081, 25113, 
    27680, 27282, 29880, 30467, 30842, 30818, 30649, 29328, 24201, 22443, 
    18785, 15477, 13887, 9091, 3336, -1361, -6115, -8973, -12418, -16292, 
    -19636, -23516, -25288, -27616, -28644, -31586, -30973, -29900, -29818, 
    -27643, -24880, -22498, -20093, -16757, -12320, -7965, -3673, -146, 3174, 
    8067, 13027, 16383, 20189, 23097, 26618, 29531, 29955, 30091, 31848, 
    29599, 29548, 28523, 25569, 23563, 20385, 16685, 11315, 8206, 5259, 21, 
    -3400, -9612, -14083, -15503, -20813, -23085, -24926, -27126, -30586, 
    -30444, -31070, -29821, -30583, -28571, -25960, -22395, -18338, -17942, 
    -14082, -7404, -3465, 608, 5058, 7505, 13433, 15999, 20278, 22102, 25101, 
    28074, 28847, 30563, 30706, 31392, 30771, 27181, 26721, 23296, 20016, 
    16680, 13945, 8615, 5368, -277, -2745, -8683, -12845, -17630, -19847, 
    -23475, -24433, -29158, -29905, -30100, -30497, -30243, -30162, -29083, 
    -25820, -23546, -21326, -16092, -13951, -8716, -3979, 415, 3430, 8943, 
    13845, 14983, 20036, 21738, 24763, 27422, 30058, 30388, 31747, 30966, 
    30718, 26909, 25890, 22766, 19799, 17086, 13383, 9135, 5395, 691, -3672, 
    -8148, -13004, -16651, -20542, -23473, -25683, -28170, -29883, -31422, 
    -31416, -31136, -29903, -29142, -27187, -24305, -20743, -16488, -13088, 
    -10751, -6223, -1559, 3248, 7525, 10676, 15578, 20066, 23610, 24740, 
    26182, 29553, 29203, 30956, 30636, 28672, 27143, 26073, 24195, 21087, 
    17472, 12786, 10508, 6036, 1469, -3394, -7689, -12862, -15678, -18590, 
    -21646, -25766, -29105, -28126, -29856, -30980, -31187, -30355, -28281, 
    -26117, -24066, -20599, -17827, -14502, -10378, -6066, -1619, 2531, 6791, 
    12755, 16161, 18141, 22272, 25892, 27686, 29915, 30875, 30396, 30033, 
    31745, 28754, 26602, 25043, 22106, 17481, 13091, 10038, 5094, 2738, 
    -2333, -7660, -11923, -14138, -18240, -22730, -25685, -26314, -30827, 
    -31034, -31476, -31491, -29482, -27125, -25502, -24535, -23321, -17101, 
    -14693, -9099, -7031, -1811, 3107, 6736, 11531, 15067, 18510, 22929, 
    24781, 28779, 28769, 30588, 30740, 30895, 30170, 29375, 27848, 23277, 
    20958, 18480, 14308, 9291, 6788, 3616, -2341, -6702, -10829, -16795, 
    -18394, -21135, -25877, -25696, -28628, -29914, -29552, -30023, -31101, 
    -29367, -27709, -25633, -20187, -18889, -13293, -10420, -6376, -3142, 
    3413, 6908, 11011, 13951, 17387, 21707, 24704, 27543, 30036, 30594, 
    29175, 31705, 28471, 29924, 27633, 24163, 21998, 18924, 16320, 11642, 
    5305, 1364, -1519, -7628, -9820, -14126, -18586, -21888, -24218, -26534, 
    -29346, -29303, -29256, -30175, -30463, -28703, -27712, -23854, -21140, 
    -19855, -15434, -11875, -6911, -1279, 509, 5162, 10613, 12882, 19079, 
    22366, 24819, 26659, 29423, 30193, 30395, 29561, 29510, 28963, 26915, 
    25129, 22319, 18890, 15326, 11531, 8684, 2286, -3132, -4343, -9638, 
    -13704, -17704, -21252, -24190, -27116, -28993, -29678, -30312, -32295, 
    -29494, -29281, -28066, -24695, -22887, -18980, -15138, -11149, -7949, 
    -4058, 1326, 5621, 10801, 12729, 16608, 21446, 24363, 26550, 28592, 
    30803, 31864, 31323, 31641, 28245, 27174, 25455, 21051, 20311, 15314, 
    10446, 7793, 2965, 252, -4236, -10946, -13763, -19005, -20855, -24129, 
    -26980, -29908, -31201, -32396, -29612, -31116, -29709, -27177, -24477, 
    -22181, -20549, -14198, -10745, -6432, -2892, 2342, 6736, 10516, 15114, 
    16581, 20115, 24417, 27772, 27472, 28860, 29968, 29266, 31224, 29999, 
    27336, 25739, 22357, 18882, 15774, 11059, 7025, 2131, -603, -4432, -8449, 
    -14174, -16209, -20930, -24424, -27672, -28305, -30347, -30226, -29902, 
    -30198, -28939, -29431, -25699, -23766, -20080, -16270, -13397, -8277, 
    -4858, -142, 4387, 7959, 14105, 16906, 20003, 23379, 25135, 27724, 29625, 
    29563, 30679, 30463, 29829, 27986, 26867, 22385, 18859, 16368, 12807, 
    9788, 4248, 771, -3480, -8771, -14309, -16963, -19886, -23563, -26258, 
    -27544, -30636, -30471, -30991, -30233, -28745, -26652, -27613, -23534, 
    -19939, -17559, -14116, -9110, -3122, -207, 4237, 8695, 12691, 17078, 
    18527, 23584, 26603, 29903, 29399, 29715, 30608, 31178, 30527, 27304, 
    26584, 24899, 20118, 17254, 12797, 7407, 3202, 161, -3846, -8046, -11375, 
    -18254, -20168, -22429, -26757, -28597, -30549, -30311, -29793, -31358, 
    -28889, -28631, -26995, -23272, -20141, -17450, -12134, -8527, -4188, 
    -227, 4437, 7996, 11571, 16311, 19311, 21920, 25081, 28194, 30301, 30341, 
    30750, 30017, 28175, 28191, 27211, 23370, 20312, 16987, 12107, 8360, 
    4362, 468, -3196, -6887, -12865, -15305, -19089, -23253, -26851, -26798, 
    -29384, -29497, -29891, -30528, -30591, -28076, -27170, -24510, -21313, 
    -15978, -13612, -9278, -5103, -88, 3103, 7670, 12970, 15062, 18763, 
    23259, 26044, 27982, 29295, 28637, 30678, 30672, 28861, 29350, 27344, 
    25351, 20398, 17679, 13777, 8704, 5340, 1826, -3687, -6449, -10598, 
    -14865, -19549, -23214, -26410, -28540, -29744, -31255, -30151, -29939, 
    -30735, -28228, -26174, -24802, -22315, -17659, -13485, -11127, -6139, 
    -2468, 3387, 7155, 12364, 16095, 19390, 22311, 24189, 25997, 30033, 
    28630, 30216, 30366, 29928, 29503, 26666, 23889, 19986, 18046, 14511, 
    10626, 5411, 953, -2287, -6864, -11619, -14001, -19887, -22150, -24890, 
    -27633, -28831, -30059, -31341, -30386, -30164, -28205, -26744, -24215, 
    -22224, -18289, -14680, -11016, -6471, -1094, 2479, 5787, 11051, 15307, 
    19325, 21921, 24267, 26917, 28974, 30800, 31330, 31085, 29891, 29159, 
    26386, 24800, 21910, 17602, 15319, 11332, 6700, 1665, -2974, -6218, 
    -11282, -16293, -17810, -22955, -25001, -26844, -27728, -29049, -29612, 
    -30961, -30833, -30222, -27378, -24511, -22810, -17494, -14810, -9550, 
    -6153, -2536, 1541, 6504, 10756, 15423, 18818, 21732, 24533, 26435, 
    28215, 30961, 29846, 30927, 30088, 29963, 27250, 24886, 20756, 18438, 
    16122, 10910, 7078, 1600, -2192, -5805, -9569, -13545, -18698, -20822, 
    -25236, -26897, -29492, -30719, -31845, -31144, -31464, -29787, -27485, 
    -24953, -21779, -18184, -14725, -10187, -6666, -1832, 1526, 5489, 9716, 
    13922, 18506, 21894, 22999, 26890, 28398, 30275, 29949, 30480, 30026, 
    29670, 27074, 26590, 22014, 18746, 13776, 11904, 6193, 3710, -2032, 
    -6180, -10412, -12668, -17191, -22115, -22580, -27601, -28038, -30043, 
    -30684, -31469, -29540, -29727, -27182, -26356, -22056, -18683, -15875, 
    -13096, -8031, -1364, 449, 6578, 9902, 13793, 17170, 20480, 23232, 25183, 
    28898, 29266, 31048, 30961, 31945, 28298, 27487, 24949, 21871, 19446, 
    15129, 10663, 7129, 3944, -552, -5602, -9827, -14470, -18115, -20968, 
    -23494, -27545, -28579, -31405, -30559, -30772, -29605, -29407, -27595, 
    -25907, -22106, -18991, -16233, -11435, -8385, -3009, -82, 4081, 10190, 
    12448, 16802, 20116, 22159, 27441, 27550, 31049, 29650, 31860, 31296, 
    29898, 28553, 27114, 23436, 18674, 16584, 11486, 7851, 3710, -2021, 
    -4838, -9817, -14313, -17111, -21075, -24279, -26193, -29702, -31030, 
    -31475, -31701, -30695, -30024, -27731, -24134, -22293, -19713, -16417, 
    -11432, -7899, -4662, 1431, 3997, 8730, 13454, 15503, 20523, 22649, 
    26255, 27640, 28542, 30506, 30050, 30062, 30245, 28711, 24706, 23336, 
    19397, 18130, 13118, 7727, 4373, -457, -4650, -7467, -12970, -16701, 
    -19098, -23024, -24553, -29236, -30997, -30743, -29225, -29761, -28676, 
    -27696, -26537, -22023, -19576, -16566, -12153, -7378, -5012, 270, 3925, 
    8741, 12513, 17405, 20296, 22300, 26009, 26928, 30031, 30044, 32000, 
    30153, 29301, 28155, 25995, 25035, 19034, 17472, 14147, 7715, 3192, 1385, 
    -3773, -9835, -12409, -15640, -19649, -22326, -26303, -26737, -28480, 
    -31047, -30717, -29504, -30439, -28479, -26257, -25120, -21172, -17618, 
    -12961, -9271, -4937, 256, 3595, 8255, 12123, 16836, 20141, 23104, 25002, 
    27560, 29868, 30398, 30539, 30201, 29598, 27792, 25341, 24450, 19987, 
    17279, 12122, 8144, 4339, -241, -5155, -8464, -12081, -16267, -19665, 
    -22779, -25819, -26441, -30721, -31504, -31836, -29182, -29839, -28373, 
    -26106, -22392, -21647, -17197, -13664, -11400, -5470, -1100, 3223, 8824, 
    12420, 16973, 19787, 23147, 24244, 28014, 29190, 29673, 29698, 31584, 
    28280, 27746, 26600, 24236, 22174, 18331, 13833, 9865, 4142, 1015, -3257, 
    -6899, -11523, -14820, -20481, -22775, -25823, -29054, -29706, -28920, 
    -29806, -31468, -29716, -29574, -28054, -23252, -21378, -17709, -13251, 
    -8953, -4330, -2686, 3371, 6235, 11247, 14984, 20249, 21417, 26093, 
    28151, 30889, 29160, 30232, 32318, 30073, 29265, 27159, 24281, 22871, 
    18010, 15939, 9129, 5017, 3133, -2918, -7844, -11480, -15576, -19008, 
    -22676, -26390, -27906, -29771, -31201, -31352, -30325, -29484, -29716, 
    -27069, -25637, -21471, -17381, -12952, -10565, -6539, -81, 2322, 6024, 
    11530, 13884, 19783, 22139, 24605, 26007, 28274, 30388, 30153, 30148, 
    28644, 30294, 26774, 25289, 21887, 18038, 14292, 9416, 5583, 1968, -1790, 
    -6652, -11657, -14373, -16897, -21703, -24133, -26982, -29069, -30427, 
    -30047, -30523, -31379, -29455, -26838, -23350, -21728, -17344, -13986, 
    -10174, -6359, -1872, 2739, 7379, 10654, 14471, 17110, 23060, 24564, 
    25771, 28230, 29738, 30664, 31039, 30247, 30289, 26172, 24124, 22375, 
    18112, 14691, 11455, 5841, 2876, -2408, -6681, -10875, -13727, -18498, 
    -21140, -23547, -28326, -28719, -30840, -30753, -30644, -29694, -28868, 
    -26817, -25529, -21069, -19513, -15786, -11855, -6655, -3708, 2256, 6029, 
    10747, 14557, 18054, 22693, 25028, 25838, 27233, 30048, 29901, 29903, 
    30228, 28716, 27133, 26154, 23361, 18773, 14014, 12433, 7968, 2690, 
    -1427, -5968, -9684, -15088, -17691, -22199, -25516, -27716, -28856, 
    -30668, -29888, -31891, -31584, -30172, -27247, -24153, -22313, -19083, 
    -14696, -10423, -5705, -3654, 3026, 6329, 9040, 13530, 18366, 21248, 
    25732, 27739, 29658, 30374, 29817, 31712, 31818, 28891, 26249, 26014, 
    23482, 17959, 15835, 10575, 6935, 2307, -719, -5786, -9535, -13559, 
    -16255, -22412, -24081, -26375, -29025, -29702, -29173, -31813, -29795, 
    -29267, -28849, -24200, -21893, -18921, -14848, -13355, -9755, -4417, 
    1353, 5682, 11059, 12557, 17175, 21075, 23277, 25178, 26710, 28846, 
    30908, 29338, 31373, 27730, 27639, 24807, 24208, 20676, 14483, 13105, 
    7817, 5180, 476, -4124, -8593, -12505, -17483, -20294, -23120, -25668, 
    -29090, -29585, -30484, -30188, -30281, -31086, -27152, -25717, -23392, 
    -19155, -16165, -12639, -7183, -4409, 168, 3708, 8349, 12357, 16319, 
    20775, 24315, 25601, 29302, 28960, 30360, 31444, 30369, 30287, 27944, 
    25450, 22875, 20976, 17442, 12652, 7660, 3672, -691, -3273, -7727, 
    -11457, -16391, -20499, -22431, -26176, -28662, -30692, -31131, -31484, 
    -29767, -28503, -28693, -25819, -24341, -20870, -16475, -13495, -9244, 
    -4830, -390, 3186, 10133, 14352, 17267, 20507, 23287, 26580, 28526, 
    29789, 29395, 31589, 29402, 30744, 28093, 25570, 22728, 20381, 16783, 
    13662, 9876, 3796, 84, -4268, -9224, -11986, -15670, -20006, -23727, 
    -25315, -27032, -29523, -29388, -30342, -30747, -30317, -28840, -26983, 
    -22948, -20564, -16061, -13050, -9677, -3648, -1182, 4655, 8410, 11658, 
    15616, 19033, 22402, 26714, 27561, 29363, 30439, 31256, 31413, 27933, 
    28979, 27432, 23028, 20536, 18383, 11723, 9033, 4749, 1230, -3792, -8197, 
    -12401, -16863, -20081, -23516, -25149, -27466, -30136, -30488, -30562, 
    -29740, -29478, -28955, -26404, -23376, -20642, -16833, -14450, -8896, 
    -5599, -844, 2477, 8635, 10638, 16460, 19977, 22019, 24356, 26443, 29469, 
    29917, 31305, 30840, 30619, 28631, 25982, 24232, 21233, 18195, 13191, 
    10105, 5198, 1186, -3202, -7834, -12668, -15929, -19262, -23960, -25154, 
    -26430, -28918, -29778, -31549, -29367, -30092, -28799, -27228, -23988, 
    -20951, -18153, -14305, -9568, -5473, -798, 3761, 7447, 11191, 14313, 
    20125, 22159, 25587, 27719, 28316, 29979, 30723, 29486, 29280, 28613, 
    27508, 24918, 21812, 16897, 13516, 10340, 7104, 1892, -2498, -5947, 
    -12003, -14815, -18522, -22829, -25179, -26644, -30891, -31353, -30783, 
    -29522, -28277, -29121, -26923, -23603, -22484, -18921, -15821, -10694, 
    -4924, -1063, 3991, 6834, 9867, 15281, 20558, 21627, 24500, 26092, 28270, 
    30322, 30691, 30510, 29591, 28253, 27006, 25979, 22098, 18511, 13967, 
    9771, 5493, 2058, -2568, -7287, -10879, -16037, -19120, -21452, -24999, 
    -27288, -27646, -30250, -30670, -30705, -30432, -28907, -25592, -24327, 
    -21819, -18242, -13320, -11902, -6433, -2358, 3049, 8379, 10252, 14068, 
    19795, 22443, 25740, 26699, 27543, 31177, 30424, 30018, 30988, 28136, 
    27804, 24631, 20891, 18826, 14540, 9609, 6857, 3558, -2056, -5250, -9606, 
    -13865, -17056, -21478, -26313, -26351, -30201, -30099, -30329, -30053, 
    -31166, -28958, -26988, -25163, -21630, -18500, -16086, -10468, -5838, 
    -2874, 1260, 7018, 9581, 15188, 18129, 22159, 23806, 27960, 28900, 29989, 
    30274, 31458, 30040, 27255, 27682, 25426, 21749, 20524, 16099, 10109, 
    6281, 3732, -2525, -4886, -9357, -15136, -17458, -20188, -23548, -25412, 
    -28466, -30172, -31469, -31471, -30605, -30104, -28353, -25829, -24159, 
    -19207, -16343, -12401, -6696, -3281, 809, 5700, 10098, 14806, 17573, 
    21214, 24638, 27223, 28431, 31211, 30477, 30391, 31078, 29408, 25859, 
    25501, 22750, 18687, 16196, 11879, 6832, 2749, -483, -5562, -9767, 
    -13907, -16402, -19888, -24319, -27143, -28941, -28474, -31135, -30976, 
    -30780, -29973, -26305, -25209, -21311, -19131, -16017, -11007, -7957, 
    -2546, 839, 6221, 10510, 13227, 17455, 20103, 23942, 25947, 29116, 30336, 
    29392, 31826, 31094, 29666, 27567, 24615, 23234, 18847, 16075, 12790, 
    7362, 4656, -1270, -5513, -8999, -13256, -18208, -20304, -23724, -27448, 
    -28778, -31133, -30520, -31686, -30583, -29963, -27072, -26149, -24087, 
    -18867, -17082, -12543, -9574, -3922, -164, 5416, 8615, 13251, 17268, 
    19924, 23907, 26627, 28628, 30503, 31012, 32071, 31358, 29511, 26759, 
    26931, 22310, 19576, 17471, 12186, 9271, 4331, -402, -4916, -10087, 
    -14506, -16290, -21184, -23816, -25603, -29172, -29244, -30615, -32086, 
    -30905, -31038, -28087, -25171, -24496, -20051, -16237, -11861, -8928, 
    -3929, 1410, 4468, 7329, 12240, 17128, 20531, 22229, 25323, 28033, 29450, 
    30560, 31190, 31048, 28172, 29146, 26757, 22696, 21787, 16967, 14599, 
    9164, 3112, -377, -3637, -8368, -10835, -17260, -19544, -24422, -25140, 
    -27896, -28687, -30328, -30320, -30560, -29995, -29199, -26008, -24010, 
    -21145, -15666, -13226, -9358, -5172, 162, 4134, 8565, 13133, 15780, 
    20107, 23971, 25121, 28348, 29311, 30734, 29447, 30134, 29013, 30033, 
    24894, 22407, 20065, 17376, 13548, 10484, 4504, 1184, -3328, -8511, 
    -12469, -14966, -19067, -24167, -25524, -27832, -29868, -30894, -30917, 
    -32395, -29846, -26894, -26402, -23674, -21499, -18686, -12738, -9772, 
    -6288, 98, 3338, 8578, 11633, 15890, 20103, 23784, 25736, 28551, 28427, 
    30240, 31019, 31744, 29886, 26671, 25075, 23465, 20724, 19190, 13733, 
    9349, 5492, 1525, -2265, -9042, -12109, -15579, -18611, -21963, -24002, 
    -28519, -29360, -31066, -30629, -30465, -31245, -28432, -26780, -24366, 
    -21994, -18149, -12359, -10278, -6010, -2417, 1219, 6416, 12075, 15262, 
    18031, 20669, 24341, 28931, 30169, 29337, 31684, 30477, 28565, 30123, 
    27955, 22617, 20502, 17376, 13847, 11057, 6843, 1707, -2307, -8675, 
    -11085, -14542, -18685, -22899, -23807, -27905, -29781, -30557, -30015, 
    -30729, -30207, -29536, -25801, -23711, -22301, -18351, -14966, -10523, 
    -5766, -1217, 2535, 6067, 11734, 15050, 19199, 22569, 25582, 28129, 
    27954, 30997, 31289, 31284, 29609, 28025, 26589, 24891, 21699, 19062, 
    14189, 11062, 7331, 3395, -2748, -7352, -11029, -14845, -18721, -23216, 
    -23382, -26514, -28782, -30090, -29961, -31418, -29952, -29505, -26110, 
    -23147, -22500, -18543, -16023, -12418, -6917, -2237, 1224, 6441, 11794, 
    15822, 18801, 23224, 23937, 27475, 28642, 29942, 30179, 30983, 29388, 
    28545, 26659, 25582, 21566, 17988, 16018, 12449, 7230, 3231, -2432, 
    -5800, -9906, -14678, -18670, -21039, -25535, -28231, -29913, -29985, 
    -30631, -31090, -29889, -27371, -26980, -25801, -23255, -20284, -15167, 
    -9729, -8509, -3172, 399, 6440, 10413, 13149, 18526, 21321, 24431, 27042, 
    28806, 30318, 30972, 30340, 29755, 29936, 27359, 24770, 22578, 18991, 
    16520, 9824, 7409, 2267, -398, -5563, -10210, -15008, -17251, -21778, 
    -23765, -25993, -28694, -29231, -30918, -31359, -28704, -30205, -27143, 
    -25116, -22573, -19697, -14669, -11214, -7430, -2727, 764, 5634, 10801, 
    14071, 17394, 21678, 24010, 25121, 27432, 29865, 30138, 32093, 29870, 
    28535, 27066, 25826, 22800, 19261, 16899, 11646, 7950, 3232, -915, -5664, 
    -8171, -14036, -16472, -20677, -24045, -26889, -28327, -30873, -30289, 
    -30369, -29862, -28862, -28125, -26990, -22777, -19675, -14501, -11748, 
    -6850, -4568, 207, 4462, 9391, 12273, 15722, 20365, 23520, 24980, 28437, 
    28860, 30455, 30700, 29185, 30120, 28506, 25651, 23251, 18250, 16384, 
    11497, 8231, 3462, 446, -5548, -8781, -13809, -18898, -18885, -24341, 
    -27152, -28693, -28468, -31163, -32332, -30125, -28652, -28327, -25787, 
    -22408, -19219, -15667, -12534, -7623, -4248, 673, 5883, 8794, 13317, 
    16653, 20447, 23651, 25582, 29076, 28864, 31623, 30751, 29944, 29709, 
    27906, 25792, 23112, 21272, 15465, 13312, 8453, 2853, -841, -4660, -8183, 
    -13693, -17603, -18661, -23764, -24618, -27486, -29914, -30070, -30300, 
    -29915, -27996, -29285, -27452, -24174, -18851, -16229, -12652, -7984, 
    -5758, -989, 4884, 8887, 12710, 15546, 21992, 24288, 25425, 29248, 29015, 
    30088, 29928, 31447, 29727, 26978, 27556, 24182, 21238, 16688, 13347, 
    8746, 3581, 507, -4420, -7728, -12128, -15769, -19028, -24446, -25796, 
    -27677, -29344, -30707, -30286, -30564, -30612, -28761, -26480, -21991, 
    -20645, -17562, -14688, -9540, -5562, -1292, 4720, 7127, 12402, 16094, 
    19341, 23370, 25905, 26719, 29644, 30049, 30604, 31567, 28551, 28849, 
    26605, 25125, 20718, 17214, 12777, 9733, 5438, 985, -4874, -9005, -10804, 
    -15697, -19715, -22232, -24312, -27953, -28031, -30247, -29189, -30118, 
    -29057, -27989, -26130, -23506, -20981, -17459, -13355, -10150, -6227, 
    -237, 3489, 8110, 11490, 14834, 19290, 23036, 24465, 27400, 29549, 28723, 
    31555, 29742, 29926, 27709, 26527, 22997, 22419, 16414, 14238, 8711, 
    4585, 2180, -3766, -7473, -11546, -16039, -19748, -21163, -24503, -27261, 
    -28635, -31418, -32086, -31265, -29543, -29637, -28012, -22565, -21291, 
    -17356, -13774, -10895, -5297, -2200, 3586, 7361, 12013, 16299, 19898, 
    23635, 26691, 27930, 28617, 30262, 30822, 31433, 28606, 29035, 26626, 
    24020, 23065, 19109, 14019, 10919, 5383, 924, -3871, -7919, -11743, 
    -15374, -18453, -21280, -24715, -25951, -29884, -29791, -31151, -30337, 
    -30603, -28496, -26072, -24646, -21785, -18365, -13286, -9927, -6038, 
    -1779, 3129, 5753, 10645, 14624, 17994, 23069, 24897, 26921, 29977, 
    30036, 30032, 30701, 30451, 30489, 26760, 24700, 22345, 18880, 15127, 
    11131, 6522, 2222, -1383, -5438, -9984, -14319, -18928, -22414, -24376, 
    -27395, -29541, -28767, -31690, -32052, -29458, -29881, -26310, -24191, 
    -21491, -17797, -14863, -10414, -7268, -3146, 2490, 5923, 11278, 15493, 
    18092, 21483, 24796, 26017, 28041, 29539, 30480, 31179, 31259, 27572, 
    25812, 23568, 21652, 17827, 16548, 11719, 6074, 2579, -1989, -7708, 
    -10225, -14236, -18338, -22660, -25762, -26495, -27849, -29779, -30075, 
    -31695, -28859, -27682, -26175, -25182, -20736, -17832, -15739, -11467, 
    -7298, -2972, 2545, 6293, 11866, 12885, 17553, 21585, 25048, 26567, 
    27169, 31350, 30642, 31572, 30082, 30460, 27499, 24658, 22329, 18620, 
    15649, 11068, 8002, 1974, -2455, -5274, -10919, -12544, -18197, -21218, 
    -24551, -25883, -27579, -28825, -31052, -30847, -30823, -29556, -27486, 
    -25271, -22160, -19121, -15954, -11229, -8345, -2972, 2437, 6235, 8257, 
    13937, 18422, 22650, 25476, 27746, 26803, 31686, 29046, 32047, 30389, 
    29837, 26212, 24945, 23448, 18026, 15885, 10940, 6806, 1746, -1847, 
    -4515, -10146, -14055, -17584, -21717, -22268, -25400, -28726, -29015, 
    -30518, -30246, -30840, -30121, -26523, -25661, -22504, -18783, -15726, 
    -12388, -7842, -3520, 749, 4939, 9216, 12772, 17436, 19871, 23138, 26157, 
    29436, 29947, 30549, 30416, 29090, 28305, 27401, 24637, 22970, 19362, 
    16566, 11689, 6681, 2008, -1576, -4723, -9313, -13659, -16609, -20476, 
    -23654, -25663, -27598, -28355, -31863, -30947, -30071, -29359, -25968, 
    -25942, -22370, -20511, -17207, -12625, -7697, -3581, 76, 5618, 10140, 
    12456, 16905, 20696, 23448, 26596, 28666, 30016, 30738, 31463, 30340, 
    30492, 28558, 25286, 24269, 19223, 15713, 12829, 7131, 2439, -97, -4843, 
    -9546, -12513, -16449, -20519, -22867, -24349, -28008, -29380, -29723, 
    -32043, -30538, -28153, -27914, -25211, -24815, -19936, -16983, -13033, 
    -8522, -4989, -553, 5613, 9047, 11449, 15675, 21847, 23617, 27051, 27859, 
    29388, 30950, 30478, 29703, 28803, 26968, 27458, 24655, 18965, 16346, 
    13094, 9479, 4557, 238, -4841, -8597, -13360, -17934, -18871, -23204, 
    -26559, -29689, -29862, -29229, -30838, -28838, -28215, -27336, -25655, 
    -22751, -19604, -16581, -11496, -10161, -3645, -138, 5481, 6529, 12933, 
    15168, 18854, 22802, 26576, 27216, 29221, 29479, 31322, 30866, 29494, 
    28873, 25935, 22870, 20172, 16701, 13933, 7355, 3775, 1413, -3695, -7906, 
    -12428, -16743, -19592, -22328, -26527, -28805, -29515, -30743, -31273, 
    -29815, -30553, -29411, -24936, -25733, -21135, -15934, -14015, -10765, 
    -6431, -2307, 3936, 7167, 12236, 17131, 19013, 22078, 24859, 25932, 
    30279, 29788, 30952, 30776, 29654, 27088, 25830, 24140, 21568, 17492, 
    14721, 9726, 4293, 1892, -3685, -6599, -11268, -14618, -18163, -21297, 
    -24787, -26752, -29454, -30628, -31465, -31527, -30543, -28402, -26568, 
    -25000, -21731, -19044, -13518, -8294, -5879, -1029, 4037, 6848, 11014, 
    15108, 18864, 21944, 25224, 25779, 28380, 30750, 30677, 29556, 28714, 
    28658, 27108, 25314, 21283, 18933, 15264, 9025, 6297, 1957, -1578, -7594, 
    -11561, -15523, -19376, -22435, -24460, -27771, -28216, -30290, -31153, 
    -30155, -29011, -29824, -25498, -25124, -20927, -16753, -15754, -12219, 
    -5841, -1796, 3265, 6816, 11492, 14538, 18126, 21313, 25477, 26451, 
    28820, 30001, 31364, 32156, 29729, 27583, 28079, 24772, 22520, 17306, 
    13924, 10983, 6287, 2662, -1662, -6711, -12386, -14517, -18811, -21837, 
    -24129, -27333, -29956, -30147, -29929, -31225, -28294, -28382, -27234, 
    -25570, -21939, -18624, -15178, -11024, -6839, -2472, 2618, 7790, 10212, 
    15480, 17569, 21847, 25746, 26244, 29193, 30704, 32070, 30093, 30468, 
    29574, 26429, 24087, 21234, 18509, 14995, 11519, 6618, 2402, -2076, 
    -7552, -11832, -14314, -17802, -21801, -24807, -28221, -27842, -29915, 
    -29832, -30219, -30681, -29149, -26624, -26108, -21902, -19222, -14075, 
    -12083, -7448, -3801, 1573, 5548, 10760, 14260, 18380, 22067, 24198, 
    28091, 28944, 30309, 32050, 29341, 29562, 29632, 27565, 25301, 22487, 
    20037, 16141, 11976, 7077, 2695, -2979, -5741, -9121, -15134, -19494, 
    -22384, -23793, -27934, -28766, -29385, -30657, -32537, -31558, -28419, 
    -27945, -24899, -21981, -19279, -14939, -10131, -8101, -2867, 340, 5460, 
    10712, 14344, 17119, 22661, 23902, 25665, 28713, 30254, 30357, 31088, 
    30230, 28065, 27197, 25784, 23277, 17743, 16731, 12540, 7629, 3761, 
    -1636, -6709, -9133, -12794, -17574, -19251, -24547, -26034, -27995, 
    -29686, -29628, -31196, -30485, -28086, -26616, -26808, -22444, -20178, 
    -15303, -12575, -7625, -4583, 1654, 5435, 9485, 13444, 17714, 21583, 
    23686, 25920, 29200, 29572, 30761, 31455, 29897, 28478, 28416, 26201, 
    24034, 19874, 15973, 12904, 8742, 3509, 386, -5090, -8012, -12856, 
    -16618, -21455, -23750, -26121, -29029, -31135, -31304, -31658, -31141, 
    -29136, -28301, -24982, -22088, -20814, -14705, -12803, -8003, -4472, 
    398, 5587, 9873, 13415, 15739, 20311, 24036, 26465, 27596, 29730, 30671, 
    32380, 30727, 29480, 29145, 26335, 22128, 19827, 16388, 12486, 9270, 
    3797, 1179, -5418, -8379, -12202, -15970, -21122, -24096, -24720, -28928, 
    -29648, -30714, -30488, -30064, -29503, -27708, -25681, -24006, -18873, 
    -16316, -12600, -8004, -4997, -47, 3829, 7433, 12188, 15246, 19927, 
    22803, 25466, 27132, 29220, 30912, 30640, 30219, 29482, 28527, 26264, 
    22401, 20868, 15145, 12057, 7745, 4568, 16, -4439, -9801, -12196, -15498, 
    -19968, -22312, -25882, -29432, -29173, -30061, -31445, -31137, -30178, 
    -26726, -24997, -24335, -20340, -17393, -11983, -8922, -5155, 857, 4566, 
    8537, 10791, 17931, 20579, 22076, 25258, 28650, 29357, 29491, 31653, 
    28816, 29099, 28941, 25094, 23874, 19590, 16277, 12990, 9013, 5262, 367, 
    -3047, -9421, -12900, -16010, -19393, -22938, -25216, -29101, -29341, 
    -30625, -30942, -29512, -30167, -27796, -26875, -22861, -20362, -15742, 
    -13118, -11106, -4174, -1299, 3582, 7127, 12063, 15646, 18522, 22921, 
    25726, 27530, 27914, 30418, 31695, 31194, 31091, 27820, 26987, 23474, 
    21873, 17161, 14049, 9006, 3789, 710, -3194, -7011, -11673, -14315, 
    -18820, -21473, -25468, -27609, -29161, -29036, -29270, -30936, -29694, 
    -27754, -26650, -24406, -21504, -16718, -15053, -10968, -5676, -989, 
    3554, 7627, 13097, 15527, 20160, 21562, 24996, 27599, 27814, 30664, 
    30738, 29579, 30124, 28424, 25325, 23154, 21482, 17824, 13525, 10122, 
    6694, 460, -3304, -8509, -11948, -14321, -18413, -23023, -25399, -26649, 
    -29250, -29604, -30644, -30794, -29988, -29670, -28078, -23207, -21420, 
    -19279, -14698, -10138, -4864, -1369, 1849, 8503, 10775, 16005, 18688, 
    20637, 23523, 27373, 29806, 31895, 31180, 31265, 29233, 28730, 27207, 
    24854, 20907, 18089, 14785, 8907, 5786, 3445, -3910, -6778, -9195, 
    -15299, -20343, -22535, -24687, -27424, -28719, -29892, -32071, -30569, 
    -29705, -27942, -25915, -24699, -22348, -20048, -16131, -9555, -7255, 
    -2299, 3121, 6699, 10704, 15384, 16866, 22473, 23796, 27168, 28530, 
    30348, 30277, 31251, 30554, 27345, 26913, 25012, 20625, 18164, 15772, 
    10479, 6767, 3392, -2112, -5565, -10394, -16188, -18862, -22455, -25430, 
    -26678, -28381, -30127, -30203, -29474, -29575, -28878, -27805, -25034, 
    -21708, -19796, -15085, -9883, -7122, -2468, 2249, 5503, 10427, 14114, 
    18250, 21866, 25680, 26030, 27529, 29537, 31509, 29073, 31389, 28920, 
    27491, 24095, 23430, 20632, 13586, 11329, 6819, 2000, -2065, -7045, 
    -11260, -14528, -18099, -21734, -24421, -24888, -28603, -29469, -32555, 
    -30236, -29780, -28989, -28099, -24129, -22580, -18746, -16966, -10456, 
    -7203, -3910, 1796, 6356, 9311, 14606, 17888, 21715, 23203, 27868, 28523, 
    29157, 30206, 31551, 31451, 29657, 26854, 25954, 22727, 18405, 16332, 
    12785, 8673, 3169, -703, -5661, -10842, -13692, -17265, -20832, -23386, 
    -25213, -27660, -28624, -30334, -29769, -29757, -30714, -26849, -25581, 
    -23305, -20157, -14559, -10668, -7827, -3446, 1746, 4063, 8286, 12821, 
    17846, 20943, 24206, 25752, 27955, 30984, 29776, 31729, 29893, 29533, 
    26727, 25028, 21436, 19074, 15630, 12572, 6934, 2877, -1133, -5792, 
    -11109, -13087, -17773, -21419, -22244, -27100, -28332, -29020, -30086, 
    -29801, -30432, -29464, -27911, -25417, -21168, -18800, -16732, -11831, 
    -8159, -4022, 443, 4860, 9050, 12681, 16949, 21378, 24777, 24578, 28604, 
    30704, 30239, 32039, 31590, 30417, 27501, 26088, 23198, 20221, 16933, 
    13391, 8950, 3838, 673, -4912, -9193, -12441, -17178, -20703, -24482, 
    -26212, -27506, -30559, -29420, -32415, -29159, -30313, -27815, -24663, 
    -24367, -21075, -15442, -13707, -9904, -3197, 850, 3151, 8932, 12762, 
    15590, 20546, 24023, 26321, 27402, 30600, 31836, 30031, 31543, 29851, 
    28436, 26591, 23099, 21146, 16885, 13524, 8507, 4392, -438, -4442, -7664, 
    -12716, -15317, -21795, -23606, -24555, -27643, -29836, -30202, -32209, 
    -30700, -28231, -28432, -24881, -23612, -20877, -17374, -13457, -9816, 
    -5490, 795, 2499, 8861, 13926, 16182, 19508, 22818, 26473, 28018, 28477, 
    30356, 30845, 29893, 29860, 29302, 25731, 23175, 20516, 17133, 14437, 
    9619, 6369, -633, -3604, -9701, -11639, -15077, -19312, -23103, -25540, 
    -27345, -28560, -30799, -30296, -31480, -29645, -28779, -26153, -24497, 
    -22582, -17727, -12845, -10184, -4053, 208, 3039, 7246, 12820, 15326, 
    20524, 23994, 25532, 27686, 29386, 29486, 30040, 30900, 29733, 29613, 
    27200, 24102, 19356, 18199, 14300, 8960, 4951, 1453, -3476, -8939, 
    -11422, -15882, -18483, -21912, -25647, -27955, -28871, -30520, -31332, 
    -31541, -29766, -28940, -25555, -25914, -19860, -17290, -14296, -10387, 
    -5629, -1835, 2072, 6979, 10466, 14949, 20307, 22337, 26413, 26891, 
    27721, 29347, 30914, 29792, 30003, 29314, 27833, 24185, 19672, 18708, 
    14623, 10906, 5266, 2473, -3757, -7008, -11379, -15441, -19771, -21751, 
    -24072, -27058, -29131, -28676, -31270, -29471, -31210, -28653, -27763, 
    -26182, -21579, -16641, -13506, -10575, -5460, -843, 1891, 6398, 12576, 
    15451, 18378, 21305, 25522, 26879, 29647, 30090, 30249, 30196, 30087, 
    28967, 27172, 23678, 22574, 18014, 14739, 10955, 7412, 3321, -1962, 
    -8227, -10777, -13915, -19534, -21350, -25077, -26045, -29921, -29974, 
    -30917, -31456, -30089, -30278, -26997, -25755, -21849, -18624, -13960, 
    -11957, -7365, -2505, 3549, 5311, 9944, 16154, 19069, 22052, 24753, 
    28647, 30349, 29181, 30780, 31956, 31260, 27536, 26800, 24743, 22046, 
    18350, 13587, 11724, 6526, 2037, -2820, -7025, -10212, -14707, -16974, 
    -22784, -23333, -26516, -28861, -30960, -30480, -31641, -29769, -28631, 
    -28337, -24601, -21082, -17717, -14706, -11749, -7395, -1848, 2084, 4714, 
    10843, 15242, 19467, 21672, 23528, 27562, 27698, 29859, 29845, 30109, 
    29474, 29365, 27273, 25088, 23477, 18686, 14882, 11233, 5975, 3724, 
    -2894, -6933, -9592, -15985, -17731, -20861, -24750, -25226, -29531, 
    -30266, -30498, -31849, -29873, -28526, -26734, -25893, -22281, -19004, 
    -16105, -12207, -7112, -3671, 2614, 6018, 10725, 13130, 18220, 20697, 
    23994, 26900, 27678, 29666, 30886, 30879, 30954, 29335, 28426, 24720, 
    20904, 17874, 16269, 12100, 6755, 2768, -949, -5079, -10492, -12444, 
    -16536, -20152, -25006, -27012, -29477, -29624, -31244, -30695, -29352, 
    -29759, -29302, -24631, -21963, -18810, -16357, -10710, -7931, -4635, 
    985, 5895, 10041, 13384, 18057, 20381, 24038, 25668, 27948, 29885, 31131, 
    30246, 30430, 28593, 29209, 26393, 22354, 19186, 15463, 10799, 8038, 
    5379, 904, -4378, -9275, -13085, -17316, -21435, -23578, -27090, -28172, 
    -29552, -30739, -30688, -30065, -28124, -27545, -25910, -22961, -20765, 
    -16286, -13658, -7879, -3017, 854, 4250, 8229, 13448, 16139, 19473, 
    23445, 27303, 28111, 30873, 30174, 30913, 29661, 30386, 27038, 25834, 
    22225, 18879, 15917, 11718, 9207, 3076, -522, -4845, -10123, -12825, 
    -16827, -20293, -22677, -26909, -27644, -29378, -30968, -30241, -29168, 
    -28576, -28369, -26746, -22452, -21279, -16826, -11971, -8576, -3121, 
    1137, 3938, 8907, 12358, 15304, 20276, 23729, 26500, 27853, 28855, 30299, 
    29627, 32174, 29561, 28320, 26770, 23711, 19485, 16446, 13487, 7482, 
    5913, 46, -3140, -7496, -13197, -16006, -19783, -22812, -25191, -27808, 
    -29736, -31011, -29809, -31418, -27782, -29228, -27544, -23776, -20762, 
    -17020, -11518, -9071, -4650, 441, 4161, 9004, 12182, 17358, 20562, 
    23588, 24727, 28472, 29735, 30471, 29274, 31678, 30753, 29325, 26301, 
    23814, 21285, 15932, 14295, 10654, 5279, 167, -2334, -7889, -12449, 
    -16249, -18333, -22715, -25033, -28079, -27735, -30373, -30709, -28949, 
    -30209, -28742, -26544, -23494, -21722, -18291, -13464, -9907, -4193, 
    -902, 3078, 6868, 13084, 15845, 20581, 23610, 25792, 26161, 27423, 31524, 
    31066, 31087, 29131, 29634, 27001, 23142, 21032, 17514, 12814, 8471, 
    4205, 178, -2731, -9379, -11647, -16173, -19516, -21682, -25931, -27531, 
    -30139, -28896, -30548, -30096, -29703, -28079, -26442, -24175, -21531, 
    -17584, -14579, -9882, -4999, -1246, 3858, 7908, 11844, 15568, 17912, 
    20739, 25120, 28104, 28322, 31130, 30119, 29968, 29557, 29543, 27155, 
    23555, 21874, 18718, 14464, 9658, 6388, 1587, -2878, -6868, -11560, 
    -16650, -18963, -22426, -24070, -27516, -30083, -31069, -30805, -30414, 
    -30421, -28934, -27860, -24372, -21207, -18460, -13827, -11078, -7790, 
    -2421, 2708, 6474, 11523, 14683, 19325, 21737, 25734, 27296, 30636, 
    29950, 31926, 30928, 30257, 28910, 28007, 25322, 21408, 16618, 15818, 
    10397, 4731, 3014, -3015, -7573, -10050, -14643, -19001, -20789, -24759, 
    -26951, -28981, -29425, -31289, -30813, -31336, -28100, -27219, -24611, 
    -21093, -17412, -15576, -10765, -5938, -3333, 3657, 8018, 11206, 15468, 
    19104, 21136, 24610, 27394, 28464, 29524, 31430, 31918, 29339, 29442, 
    26901, 25741, 22556, 18375, 15739, 10935, 6330, 1480, -1228, -6162, 
    -9632, -13109, -18476, -21217, -24256, -27840, -27822, -29243, -30910, 
    -28995, -30656, -30039, -26734, -24161, -20897, -17884, -15802, -11286, 
    -6418, -3782, 1755, 6104, 8885, 15166, 17720, 21479, 25746, 28227, 28989, 
    29675, 30450, 31650, 30818, 28669, 25511, 25045, 22597, 20167, 16307, 
    10306, 8356, 2940, -1760, -7035, -10003, -13864, -16703, -21623, -25118, 
    -25720, -28692, -29043, -30890, -30785, -30717, -28823, -27417, -24119, 
    -22178, -19499, -15966, -12934, -6522, -2921, 740, 7507, 9664, 13830, 
    16670, 20042, 23601, 26339, 28387, 29309, 31343, 30655, 30724, 29032, 
    27835, 25993, 23076, 18686, 15474, 10297, 8474, 3150, -483, -4314, 
    -10741, -12893, -15931, -22055, -22891, -25865, -28964, -30707, -30662, 
    -30861, -29782, -29430, -26461, -25136, -23521, -19455, -16035, -13160, 
    -7994, -4044, 1114, 4345, 10168, 13921, 16753, 22270, 22968, 24799, 
    28062, 30627, 30126, 29887, 29929, 28962, 28016, 25205, 23688, 20201, 
    16746, 13097, 8916, 5002, 3, -5105, -8704, -13645, -16533, -20246, 
    -24361, -24982, -27685, -28725, -30122, -30909, -29859, -30675, -26743, 
    -25656, -23983, -20202, -17670, -12063, -8336, -4312, -647, 4036, 7733, 
    13580, 17754, 19738, 23373, 25013, 29006, 29239, 30556, 30812, 30952, 
    29020, 28748, 25368, 23443, 19988, 16989, 12625, 8428, 4265, 37, -4632, 
    -7523, -11642, -16563, -19318, -23565, -26458, -26566, -29052, -30394, 
    -31035, -31388, -28038, -27411, -26446, -23151, -20152, -16256, -14515, 
    -8138, -4375, -1692, 4357, 9098, 13007, 15741, 20114, 24393, 25816, 
    27628, 29052, 30451, 29162, 30372, 29803, 28128, 25620, 23305, 20139, 
    17067, 14527, 9260, 3993, -1525, -4630, -8193, -12628, -15696, -20407, 
    -22963, -26896, -27622, -29610, -31199, -31393, -30391, -30600, -28529, 
    -25907, -23605, -20401, -16753, -13325, -9178, -4924, -361, 2995, 7530, 
    10677, 17361, 18329, 22676, 25999, 26639, 29484, 30893, 29581, 30208, 
    29338, 29311, 26945, 24422, 21617, 16461, 12926, 10087, 5132, 1403, 
    -3057, -7890, -12324, -15743, -19692, -24015, -26512, -27380, -28466, 
    -30667, -30413, -29682, -29868, -28465, -27527, -24168, -20273, -16956, 
    -13687, -9127, -3672, -378, 2710, 8043, 12622, 16695, 19720, 22106, 
    24371, 27966, 29660, 31314, 32593, 31306, 29717, 28323, 27411, 23980, 
    19721, 17101, 15290, 10076, 4400, 1182, -1807, -7076, -11673, -15864, 
    -19466, -22118, -26366, -29059, -28619, -29504, -31274, -31132, -29342, 
    -29517, -28392, -25291, -21142, -18491, -13438, -10340, -4527, 54, 2447, 
    7428, 12107, 16361, 18011, 22099, 25174, 27108, 28247, 29943, 30785, 
    32097, 29643, 28602, 26600, 24123, 22380, 18959, 14309, 10563, 5295, 
    1678, -3220, -7346, -11150, -15988, -18363, -21474, -26114, -26113, 
    -29660, -29830, -29444, -30388, -29853, -28487, -27607, -25218, -21005, 
    -18840, -12937, -9696, -5848, -2731, 1520, 6847, 9639, 15081, 19438, 
    20960, 25542, 26465, 30570, 29588, 29777, 30704, 30097, 27816, 27647, 
    24873, 21319, 19017, 15682, 10370, 5312, 2181, -3208, -7834, -9495, 
    -14932, -17599, -23234, -26109, -27048, -27696, -30602, -31802, -29536, 
    -30961, -29109, -25495, -24397, -21204, -19395, -15717, -12249, -6686, 
    -2123, 1395, 6434, 11084, 14182, 19734, 20687, 25772, 26779, 28051, 
    31274, 31777, 32470, 31737, 27552, 27095, 24327, 21048, 19493, 14861, 
    10396, 7900, 2218, -2354, -5988, -10670, -14811, -17964, -19950, -24173, 
    -26319, -27424, -29368, -31527, -30834, -30862, -27772, -27167, -24560, 
    -21988, -18468, -14078, -10379, -7687, -2899, 1159, 5255, 9773, 15869, 
    17585, 21586, 25510, 27825, 27668, 31281, 30317, 31656, 31818, 28882, 
    25672, 26135, 22651, 18075, 16080, 11849, 6763, 3936, -1948, -4657, 
    -9945, -14288, -19281, -21624, -24509, -26228, -27481, -30319, -32086, 
    -30931, -28753, -28862, -27133, -24392, -22429, -18377, -15979, -10079, 
    -6629, -2559, 2199, 4663, 10868, 15140, 17845, 20287, 25289, 26659, 
    28473, 29363, 29756, 29638, 30341, 29417, 28846, 25133, 22665, 19048, 
    15911, 12091, 8522, 4284, -2462, -6073, -9597, -13952, -18369, -20030, 
    -23771, -26300, -27646, -29525, -28925, -31109, -29605, -29508, -27454, 
    -25412, -22783, -19421, -16045, -13022, -8079, -4248, 755, 5338, 10552, 
    14577, 16812, 20867, 25636, 27051, 28712, 30641, 31267, 31204, 31830, 
    29567, 27471, 25510, 23101, 18672, 15489, 13562, 6314, 4199, -542, -4348, 
    -9868, -12498, -17242, -21566, -24845, -24770, -28779, -29799, -30542, 
    -32481, -30009, -30071, -27218, -26662, -23430, -20161, -17611, -12713, 
    -8244, -4905, -588, 3840, 7757, 11421, 18075, 20230, 23733, 25105, 28568, 
    31469, 30011, 30672, 31071, 30556, 28464, 25453, 23503, 21179, 16692, 
    12826, 7320, 5640, -125, -3765, -8138, -13066, -16217, -20330, -23892, 
    -26408, -27381, -28827, -29489, -29705, -29752, -29574, -28055, -25743, 
    -24326, -20148, -16353, -14466, -9474, -5257, -1331, 4216, 7649, 13306, 
    16815, 20208, 23233, 25487, 28541, 30075, 29280, 30544, 29468, 28060, 
    26717, 24648, 24195, 19276, 15910, 12404, 9268, 4260, -690, -4462, -8337, 
    -12609, -17247, -20271, -23145, -25561, -28175, -29196, -30241, -30479, 
    -30282, -29392, -28459, -26131, -22974, -21183, -17483, -13094, -9988, 
    -4777, -308, 3886, 9066, 12727, 16639, 19743, 22165, 26082, 29286, 28951, 
    30876, 30528, 29540, 28686, 28964, 25434, 23185, 20844, 18695, 12725, 
    9511, 4914, 2330, -4197, -7503, -13116, -16072, -20907, -22828, -24662, 
    -27976, -29423, -28959, -30801, -31731, -29653, -28348, -27512, -24554, 
    -19330, -16450, -13842, -9620, -6817, 745, 2311, 7025, 11508, 14828, 
    20184, 23720, 25469, 27064, 30921, 30802, 31624, 30844, 30960, 28596, 
    25719, 24268, 20688, 16998, 13300, 9706, 5564, 1100, -2517, -8102, 
    -11934, -16231, -19060, -21308, -26002, -27283, -29126, -28705, -31526, 
    -30390, -30017, -28246, -28263, -23386, -20774, -17113, -13011, -10238, 
    -6757, -1031, 1467, 8344, 11778, 14332, 20383, 23191, 24104, 28153, 
    28876, 30037, 31951, 29346, 29194, 28579, 26948, 25191, 22374, 18403, 
    13390, 10316, 5992, 1212, -3479, -5548, -12016, -14406, -18874, -23533, 
    -25972, -28746, -28815, -29913, -32113, -32250, -30927, -28968, -28401, 
    -23748, -21203, -17324, -14023, -10798, -5902, -562, 1884, 5973, 12293, 
    13872, 19084, 21664, 24986, 27794, 28101, 31197, 29854, 29871, 30427, 
    28892, 26047, 24775, 22631, 18496, 14161, 10425, 6292, 2326, -3306, 
    -7336, -11282, -15417, -18982, -22730, -25289, -26404, -28240, -29081, 
    -30653, -32030, -31473, -27901, -27208, -24241, -22621, -18307, -14840, 
    -10687, -6417, -1517, 2138, 7244, 12009, 15069, 18753, 21721, 24156, 
    27505, 29210, 28908, 30422, 30887, 30090, 29035, 28242, 23727, 22475, 
    19422, 14500, 10992, 6824, 1644, -1846, -5991, -11897, -14646, -19586, 
    -21462, -26132, -28443, -29104, -31573, -30241, -31568, -29685, -29372, 
    -27162, -25990, -23427, -19032, -15302, -11568, -6757, -2395, 1704, 5279, 
    11272, 13528, 17286, 20703, 23996, 26668, 28100, 30768, 30140, 30152, 
    29943, 30041, 26380, 24947, 22307, 18768, 14130, 11751, 7685, 4690, -914, 
    -6928, -10594, -14002, -18395, -20148, -23932, -27956, -28561, -29933, 
    -30279, -29537, -29134, -28297, -26692, -25755, -22604, -18774, -15221, 
    -11974, -7315, -2511, 1398, 4338, 8610, 14709, 16698, 21007, 24687, 
    25270, 29038, 29234, 30198, 31851, 30248, 28248, 26375, 23651, 22360, 
    19371, 14297, 13487, 7690, 4471, -1193, -6275, -8924, -13093, -18657, 
    -21585, -24908, -24757, -28721, -29305, -31848, -31083, -30465, -29295, 
    -27021, -25084, -22420, -18276, -14919, -12094, -6802, -2658, 1402, 5803, 
    8696, 12373, 17742, 22375, 22957, 26158, 28077, 31355, 29885, 29900, 
    29248, 27997, 27496, 26159, 22648, 19179, 16020, 13970, 8700, 4889, 
    -1539, -4152, -8447, -14501, -16361, -20437, -23275, -26249, -29183, 
    -28657, -30007, -30758, -29279, -29368, -27854, -24417, -23875, -21361, 
    -16242, -13198, -6924, -4303, 717, 5333, 10407, 13205, 17911, 21481, 
    23925, 27114, 29053, 29680, 29229, 31589, 29908, 28594, 27414, 25413, 
    22427, 20081, 15913, 13149, 9747, 2840, 1210, -4848, -8343, -13984, 
    -17021, -20403, -23632, -25504, -27784, -29690, -31790, -30890, -31945, 
    -30216, -27413, -27372, -22600, -21505, -18228, -13681, -7803, -5370, 39, 
    3150, 7988, 14287, 16745, 20767, 23329, 26015, 27998, 31003, 29181, 
    30211, 28710, 30215, 28731, 24649, 23086, 20691, 17079, 13935, 8439, 
    4799, 291, -3859, -7408, -12545, -16055, -20785, -23048, -24501, -27712, 
    -28754, -30028, -31314, -31123, -29640, -28794, -26107, -24703, -19967, 
    -17170, -11426, -9732, -6257, -1687, 4113, 9237, 13143, 14810, 19273, 
    24246, 25543, 26199, 30208, 31330, 31606, 29206, 29615, 29438, 27481, 
    22726, 22254, 16179, 12820, 9675, 4073, -379, -2634, -8460, -11504, 
    -16558, -19076, -22754, -24813, -27587, -30605, -32061, -31241, -32293, 
    -29027, -27388, -26004, -24225, -21119, -18781, -14393, -9567, -4631, 
    453, 3698, 8475, 11452, 16080, 20499, 24164, 25713, 27252, 30260, 29360, 
    29713, 29819, 30878, 28475, 27553, 23921, 20464, 17246, 13313, 10519, 
    4194, 859, -2427, -7709, -11937, -14544, -19881, -22848, -26571, -27567, 
    -29635, -28683, -29661, -32160, -29607, -27933, -26177, -23823, -20436, 
    -17858, -12879, -9277, -4368, -662, 2664, 7650, 10510, 14290, 18377, 
    22955, 23716, 25829, 28682, 31103, 30201, 30611, 28508, 26895, 26823, 
    25391, 22057, 17780, 15554, 9891, 4895, 1682, -2527, -5972, -10698, 
    -15733, -19041, -23315, -25953, -28197, -30446, -29661, -30126, -30627, 
    -29228, -29009, -25699, -24865, -20244, -17267, -14393, -11381, -5502, 
    40, 1763, 7794, 10100, 15727, 19713, 20648, 24927, 27074, 28796, 29592, 
    30877, 29827, 30808, 28543, 26172, 24879, 20112, 17703, 15193, 11903, 
    5117, 1313, -2842, -6771, -10568, -15931, -17419, -21638, -24823, -25824, 
    -30024, -29762, -30481, -29613, -29324, -27452, -26453, -25771, -20629, 
    -20206, -14943, -10972, -6338, -3044, 1837, 5794, 10736, 14887, 19469, 
    22479, 24270, 28575, 29121, 29973, 30742, 31633, 28384, 30543, 27176, 
    25419, 21329, 20026, 15366, 11255, 5505, 1695, -1157, -7152, -11416, 
    -14926, -19590, -22565, -25312, -27960, -27646, -29700, -30546, -30424, 
    -28766, -29094, -28673, -24733, -22532, -19093, -15460, -11550, -7988, 
    -2926, 1452, 6284, 11571, 14357, 18340, 22081, 24031, 27133, 27815, 
    29310, 30799, 30026, 30177, 28830, 27565, 25579, 22305, 17462, 16801, 
    11152, 6539, 4284, -586, -6480, -9649, -15302, -17507, -23094, -22949, 
    -26343, -29404, -28402, -30604, -29676, -29854, -28889, -26980, -24863, 
    -21599, -19888, -17356, -12196, -5804, -3872, 1839, 5779, 9730, 15041, 
    18447, 21129, 23971, 26959, 28582, 28908, 30488, 31146, 29037, 29047, 
    27864, 24753, 22236, 19334, 15232, 11610, 8131, 2484, -32, -5989, -9786, 
    -14004, -17376, -21257, -23571, -26891, -27969, -29373, -30323, -31239, 
    -31207, -28444, -28299, -26214, -21953, -18348, -14674, -10777, -8484, 
    -2984, -319, 5523, 8902, 13697, 16628, 21266, 22624, 26036, 28605, 28699, 
    29451, 30388, 30953, 29733, 27818, 26032, 23483, 19699, 15803, 12801, 
    8725, 4660, -660, -4940, -9334, -11845, -16515, -19573, -23834, -25668, 
    -27547, -30047, -30173, -31469, -30837, -28784, -27472, -26076, -23233, 
    -19485, -15879, -13461, -7145, -3379, 781, 4390, 9929, 13577, 16641, 
    21384, 23922, 25307, 27362, 30834, 30782, 31803, 31317, 30293, 28173, 
    26929, 23871, 19427, 17841, 12104, 7803, 4227, -1203, -3115, -9383, 
    -13795, -17599, -21208, -23266, -26204, -28474, -29128, -29376, -32124, 
    -29721, -29420, -28085, -25583, -23691, -20633, -15596, -13630, -9014, 
    -4491, 241, 4920, 8703, 11252, 15645, 18317, 21974, 25696, 27196, 29186, 
    30164, 32007, 29588, 28764, 28078, 27114, 24053, 20555, 16634, 12305, 
    7898, 3653, 398, -3753, -8234, -12264, -16200, -18838, -23230, -24211, 
    -27897, -28575, -32168, -32394, -30013, -29853, -28779, -25140, -23748, 
    -20215, -17373, -14039, -9421, -4574, 980, 3304, 7170, 14079, 17402, 
    20635, 24214, 24686, 27546, 29472, 31726, 30826, 31782, 30768, 27838, 
    25923, 22733, 22114, 18317, 13786, 8370, 4937, 1022, -3406, -9080, 
    -11688, -16017, -18995, -24418, -23930, -28675, -28302, -31189, -31136, 
    -31833, -29621, -29500, -28099, -24224, -21209, -18056, -14455, -8965, 
    -5585, -1244, 2212, 8308, 10496, 15814, 21147, 23549, 25973, 28445, 
    30025, 30401, 29800, 31126, 28801, 29221, 25243, 24990, 21302, 17370, 
    13996, 8380, 5429, -536, -3644, -8766, -12788, -15434, -20247, -22883, 
    -25762, -27389, -29140, -30250, -31529, -30499, -30776, -28503, -27471, 
    -23100, -21458, -17916, -13426, -9794, -6921, -2210, 1779, 6725, 11775, 
    14940, 19452, 22472, 25338, 25714, 29261, 30701, 30186, 30963, 31600, 
    27528, 26049, 24881, 19990, 16360, 14203, 9403, 6782, 3079, -3808, -8397, 
    -12840, -15957, -19067, -22113, -26093, -26190, -28512, -30654, -30682, 
    -31760, -31117, -27621, -28052, -24437, -21991, -19610, -14379, -10434, 
    -5472, -1306, 3659, 7930, 9702, 15452, 18737, 23679, 25176, 27090, 28804, 
    30022, 30490, 30250, 28856, 28429, 26441, 24444, 21045, 18000, 14104, 
    9472, 5910, 895, -2039, -6947, -10354, -13621, -18154, -22268, -25339, 
    -25659, -28249, -29660, -29145, -30593, -31543, -28300, -28266, -24445, 
    -22198, -19829, -14741, -10806, -7797, -2418, 2989, 8245, 9568, 14234, 
    18190, 22116, 25219, 27028, 28334, 30641, 31275, 31902, 29320, 29333, 
    28856, 25045, 22197, 18675, 13722, 10548, 6850, 2315, -2591, -5069, 
    -10222, -14232, -19653, -21552, -24847, -27905, -29291, -29150, -29259, 
    -29337, -30247, -30069, -27734, -23313, -21345, -18955, -14982, -11914, 
    -5889, -3667, 1208, 7261, 10206, 13200, 18559, 21817, 24433, 25727, 
    29682, 29817, 31716, 31196, 30389, 29415, 27411, 24044, 23046, 18954, 
    14823, 9837, 6868, 3426, -351, -7455, -9899, -14087, -16970, -20043, 
    -24257, -26515, -26879, -29236, -30104, -31064, -29096, -29494, -27557, 
    -25870, -22495, -19511, -14516, -12120, -5884, -3145, 905, 6233, 10747, 
    14029, 17471, 21173, 24372, 26292, 26802, 28860, 29557, 30923, 29961, 
    29465, 27772, 24592, 21862, 20030, 14065, 12024, 7349, 3345, -786, -4281, 
    -9426, -14242, -16167, -22026, -23257, -26169, -27598, -30143, -30687, 
    -31485, -30740, -29323, -29164, -25216, -23328, -19308, -15887, -11691, 
    -6728, -3226, 2137, 5952, 9114, 14347, 17904, 19073, 24282, 25577, 28345, 
    30051, 30287, 30757, 31980, 29288, 27669, 25503, 21601, 19658, 17044, 
    11853, 8646, 4543, 398, -5651, -10255, -11929, -17080, -21351, -23808, 
    -25785, -29996, -28708, -31712, -30772, -30423, -28708, -27777, -25745, 
    -22991, -18629, -17765, -13926, -8478, -3681, 199, 6097, 9757, 13159, 
    18662, 20564, 23472, 25923, 27224, 29186, 30593, 31723, 30104, 30433, 
    28031, 26187, 23798, 19280, 14919, 13160, 8333, 4906, -1716, -4573, 
    -8731, -13846, -16267, -20305, -25095, -25509, -27049, -29011, -30017, 
    -30336, -31557, -29438, -27784, -25802, -21651, -20170, -16204, -13190, 
    -9437, -5002, 388, 4102, 7564, 11876, 16026, 20654, 23224, 26973, 28032, 
    29010, 30444, 30423, 31731, 30709, 28085, 27216, 23900, 20951, 16934, 
    14354, 8692, 4847, 52, -4593, -9507, -11041, -16292, -19823, -22832, 
    -26380, -26624, -28206, -31016, -32014, -30716, -29052, -27458, -26124, 
    -22486, -21673, -16117, -14506, -7658, -4448, 1202, 3242, 8232, 12962, 
    14653, 18729, 24308, 26722, 27315, 28851, 31109, 30308, 30966, 29832, 
    27728, 26509, 23609, 19865, 16349, 12883, 10112, 4239, 1156, -3189, 
    -8333, -12632, -16051, -19888, -22686, -26615, -27715, -30038, -30534, 
    -29976, -30307, -30010, -27517, -27080, -22507, -20708, -15998, -14775, 
    -8760, -4217, 363, 4690, 7321, 12209, 16578, 18856, 24032, 24016, 28356, 
    29313, 30742, 31039, 31666, 28773, 27494, 26697, 23309, 21696, 18095, 
    13081, 9821, 4662, 1770, -2875, -8388, -11944, -17130, -18491, -23058, 
    -26149, -26303, -29721, -30139, -30329, -30364, -29895, -28500, -26424, 
    -23279, -21883, -16484, -15582, -8969, -6517, -1574, 2991, 7708, 11951, 
    15606, 19906, 22498, 26412, 26288, 30643, 31130, 31022, 29171, 30569, 
    28015, 26448, 23720, 20561, 17355, 14093, 9864, 5357, 1407, -3358, -5980, 
    -11455, -15113, -18836, -21700, -23888, -27576, -30370, -29672, -30390, 
    -30526, -31531, -28617, -27218, -24663, -23168, -17730, -15092, -9744, 
    -7175, -2009, 2396, 7385, 10440, 14491, 18801, 22577, 24492, 27745, 
    28684, 30366, 31348, 30423, 28978, 29002, 26876, 25123, 23147, 18448, 
    14808, 10983, 6457, 2771, -3874, -5909, -11312, -14685, -19564, -22797, 
    -25163, -27486, -28842, -29963, -31492, -30584, -30288, -29876, -26833, 
    -24852, -22129, -19199, -15999, -11496, -5279, -1435, 1646, 6223, 10181, 
    16404, 19065, 21581, 24018, 27246, 27827, 30578, 29557, 30841, 29685, 
    27755, 27706, 26101, 21816, 18292, 16369, 11840, 5912, 3433, -2159, 
    -6196, -11921, -14126, -19024, -23168, -24401, -27874, -29259, -30194, 
    -30877, -31478, -29058, -29131, -27812, -24794, -22662, -19962, -16462, 
    -11700, -7471, -3249, 1577, 4463, 10243, 13947, 17567, 21922, 25101, 
    25859, 28208, 31562, 30415, 31524, 30228, 28815, 26890, 25674, 21657, 
    18483, 14476, 11642, 7567, 2605, -1644, -6643, -9259, -13622, -18133, 
    -22275, -23286, -26787, -27880, -29652, -29657, -30990, -30410, -29070, 
    -25872, -25325, -22767, -19465, -15126, -11258, -7466, -2363, 2516, 6568, 
    9730, 12674, 17935, 21829, 24235, 27988, 27972, 31713, 30914, 30704, 
    30501, 29847, 27456, 24964, 22334, 19425, 16461, 12288, 7406, 3517, 
    -1679, -4253, -10097, -14336, -17861, -21051, -24097, -24848, -29524, 
    -29966, -29557, -31551, -31169, -28293, -27585, -24777, -24186, -18797, 
    -16636, -11618, -6874, -3491, 1210, 5132, 8826, 13318, 16320, 21140, 
    23592, 26029, 26993, 28459, 30069, 30256, 29203, 28383, 28383, 24470, 
    22780, 19802, 17078, 12247, 8438, 3648, 123, -4699, -10798, -14087, 
    -17217, -21215, -23585, -26263, -29546, -30045, -30188, -31056, -31084, 
    -29376, -27687, -26809, -21156, -20482, -16257, -12399, -7339, -4907, 
    852, 3185, 7416, 12950, 15785, 18812, 24308, 25352, 28161, 29889, 30459, 
    30069, 31435, 28103, 28536, 26693, 23457, 19450, 16547, 11616, 7905, 
    3920, -779, -5118, -9618, -13212, -17537, -21191, -22836, -26736, -29279, 
    -29275, -30660, -31659, -30327, -29934, -27730, -25374, -22685, -21006, 
    -16071, -13377, -9015, -4072, 1207, 4929, 9057, 11494, 16917, 19696, 
    23148, 26019, 28478, 28939, 31490, 31643, 30560, 29061, 28223, 26626, 
    24252, 19788, 16751, 12794, 9247, 5733, 242, -4607, -9801, -13167, 
    -15621, -18338, -24056, -25154, -26749, -31228, -29749, -29617, -31353, 
    -29698, -27965, -27136, -22833, -21298, -16407, -13081, -9515, -5713, 
    -2052, 4017, 6944, 13877, 15723, 21357, 22300, 25433, 27135, 29593, 
    29960, 31483, 32329, 31052, 28284, 27005, 21868, 19891, 16941, 14864, 
    10292, 5585, 1530, -3532, -7591, -13653, -16757, -19447, -21978, -26087, 
    -27283, -30322, -30443, -30878, -31543, -30328, -29475, -27687, -23962, 
    -20221, -17450, -13677, -11123, -7032, 953, 2460, 8303, 12238, 14621, 
    17927, 21199, 24344, 27315, 27899, 31805, 31503, 29930, 30642, 28712, 
    25876, 24253, 19850, 16712, 13294, 10365, 4725, 543, -3338, -6009, 
    -12178, -15223, -18668, -21039, -25227, -27384, -30109, -29409, -32178, 
    -31875, -29877, -28983, -25212, -23532, -20207, -17485, -12779, -9055, 
    -4804, -341, 3787, 7729, 12369, 15485, 19000, 21453, 26577, 27736, 29391, 
    30298, 31442, 31042, 29391, 28739, 26988, 23691, 21684, 18530, 14713, 
    9156, 4747, 743, -2953, -7728, -11869, -16079, -18702, -21947, -24531, 
    -28283, -28971, -30293, -31778, -30518, -31322, -27772, -26846, -24736, 
    -21711, -19365, -15141, -11315, -4905, -2147, 1814, 6695, 11078, 14126, 
    17526, 21580, 24643, 27361, 29137, 30422, 32475, 29954, 29911, 28346, 
    28350, 25796, 22024, 18070, 14272, 10917, 6575, 2440, -1493, -6492, 
    -10351, -14668, -17481, -20384, -24461, -26619, -27703, -30273, -30970, 
    -30549, -30232, -29417, -26358, -24248, -22042, -18045, -15690, -10417, 
    -7038, -2513, 1982, 7324, 9982, 13733, 17456, 22911, 25696, 27653, 28218, 
    30003, 30595, 29770, 29511, 29346, 27746, 23596, 21774, 17426, 15277, 
    10707, 7012, 2868, -1482, -6240, -10474, -15505, -16714, -21749, -24535, 
    -26993, -29804, -30431, -30227, -30635, -30115, -28297, -27063, -25779, 
    -22459, -17769, -16116, -10056, -7462, -2468, 1395, 5652, 9396, 14503, 
    18149, 21407, 24509, 26591, 28330, 29499, 28965, 31045, 28893, 30077, 
    27820, 25533, 21694, 18373, 15300, 11205, 8407, 3545, -2806, -5721, 
    -10169, -14697, -17323, -21416, -24337, -27807, -28645, -31060, -31692, 
    -29815, -29105, -29680, -28221, -24922, -22137, -18615, -16630, -11407, 
    -8017, -3754, 1393, 5798, 9502, 12496, 17725, 20364, 22635, 27710, 29791, 
    29640, 30342, 29695, 28713, 29395, 27011, 24710, 21386, 19055, 15113, 
    11882, 8414, 3556, -3019, -6917, -10246, -13969, -19233, -20431, -23075, 
    -25075, -28157, -29408, -30454, -30827, -30448, -29480, -27550, -25598, 
    -22347, -19105, -16026, -13556, -8167, -3165, 2179, 6438, 9087, 13570, 
    17889, 21273, 23737, 25381, 29077, 30547, 30951, 29934, 29524, 30135, 
    27553, 25909, 23617, 19875, 15493, 11243, 6746, 3989, -51, -6470, -9115, 
    -13779, -17796, -20344, -25460, -24492, -27101, -29552, -31633, -30318, 
    -32106, -29491, -28053, -23951, -23336, -21220, -16098, -12428, -7213, 
    -2925, 820, 4275, 9617, 11823, 18525, 19984, 24555, 24554, 27512, 28394, 
    31377, 31482, 29305, 28503, 27392, 25514, 22619, 19208, 17409, 12502, 
    7561, 4132, 700, -3134, -9623, -12758, -16199, -20468, -22804, -24844, 
    -29055, -31401, -30955, -30910, -30446, -29785, -27865, -25762, -23656, 
    -20375, -16819, -11907, -8970, -4032, 435, 4810, 9144, 12269, 15716, 
    21866, 22880, 25039, 27827, 31037, 31420, 29877, 30226, 30182, 29141, 
    25925, 22978, 20285, 15922, 13203, 7747, 4949, 166, -3773, -8902, -13463, 
    -17030, -19488, -23189, -25207, -27659, -27942, -30858, -32383, -30246, 
    -29344, -28073, -25481, -23842, -19178, -15913, -14035, -7472, -4026, 
    -542, 3473, 7330, 12207, 16768, 21462, 23092, 26698, 28286, 28447, 30287, 
    31864, 29363, 29038, 29095, 26148, 23092, 22025, 16878, 13803, 10008, 
    4298, -498, -2637, -8123, -11127, -16233, -19526, -21868, -24889, -27300, 
    -28242, -29837, -29165, -29919, -31114, -27415, -26553, -24764, -20322, 
    -16659, -13585, -10095, -4902, -145, 3174, 8103, 13199, 15849, 18606, 
    23726, 26348, 27981, 28756, 30193, 31414, 30308, 30021, 29092, 25526, 
    23363, 21057, 18176, 14108, 8226, 5265, 1232, -1932, -7207, -12051, 
    -17013, -19019, -22701, -25761, -27360, -30406, -31717, -31638, -30549, 
    -30006, -29131, -27259, -24510, -21879, -16774, -12575, -10643, -6003, 
    -695, 2255, 6227, 11186, 15832, 18496, 23990, 25860, 27757, 29646, 29757, 
    31914, 30993, 28841, 28458, 26959, 24222, 21031, 17727, 15042, 9303, 
    6521, 2186, -3735, -7784, -11656, -15057, -19678, -23126, -23462, -28352, 
    -28068, -30163, -29617, -29864, -28613, -28866, -26465, -23538, -22829, 
    -19145, -13860, -9551, -7100, -1555, 3288, 6467, 11391, 14629, 19629, 
    22011, 26161, 26767, 28148, 30512, 28980, 30430, 30020, 29044, 26067, 
    23646, 22009, 17061, 14111, 9766, 5800, 3391, -2377, -6913, -9958, 
    -15340, -18415, -21015, -26252, -26855, -29011, -30581, -30180, -30297, 
    -30096, -28305, -25977, -24473, -21263, -17779, -15239, -9325, -6129, 
    -2098, 1992, 7251, 11616, 14381, 18723, 22332, 24645, 28259, 29961, 
    29331, 31691, 29164, 29475, 28161, 27037, 23922, 22960, 18602, 13978, 
    10808, 6783, 2024, -2597, -6859, -11975, -14444, -17204, -22000, -23847, 
    -26489, -27643, -29757, -31832, -30044, -31547, -27941, -27554, -24623, 
    -20882, -17293, -15692, -12383, -7133, -3209, 912, 5247, 10346, 14615, 
    17125, 21514, 23733, 25440, 27168, 29807, 30817, 31157, 31605, 28469, 
    28871, 26248, 21842, 18580, 15018, 11419, 7986, 2293, -1230, -5895, 
    -11145, -12499, -17923, -20099, -24757, -26055, -28492, -30968, -30272, 
    -32096, -29494, -30042, -26503, -24535, -22416, -19827, -16267, -11642, 
    -7307, -3431, 1227, 5281, 8526, 14621, 18925, 22447, 23440, 25721, 27948, 
    29803, 30736, 31612, 28949, 29934, 26655, 24864, 22967, 18896, 15138, 
    12734, 8683, 2515, -517, -5158, -10121, -12016, -17651, -21548, -22192, 
    -27613, -27410, -30423, -30439, -30439, -31734, -28474, -27169, -25356, 
    -21356, -20249, -15642, -12668, -7862, -3404, -80, 4500, 8907, 13409, 
    16966, 20931, 23133, 25892, 29451, 29912, 30308, 29548, 29971, 29044, 
    27933, 24013, 22495, 19046, 16905, 12137, 8481, 3091, -477, -4316, -9056, 
    -13325, -16128, -20569, -22665, -27513, -28280, -29450, -29954, -31722, 
    -30778, -28205, -27786, -24755, -23671, -19298, -17823, -11605, -7864, 
    -2983, 47, 5194, 9066, 13073, 17187, 18984, 24777, 25686, 29040, 29787, 
    30489, 30189, 29966, 29215, 27742, 25252, 22608, 19244, 16690, 12465, 
    8378, 4265, 431, -5504, -7935, -12419, -17863, -20302, -22578, -27403, 
    -27125, -29691, -30183, -30764, -30256, -30271, -29147, -26932, -23146, 
    -19766, -16992, -12479, -8299, -4676, -839, 3827, 7577, 13865, 17824, 
    20198, 24017, 27238, 29236, 29763, 29788, 29374, 30107, 29320, 27897, 
    25965, 23803, 21104, 16646, 13204, 7426, 3421, 278, -4139, -9435, -10973, 
    -15297, -19250, -22254, -26231, -27842, -30712, -30354, -31249, -30986, 
    -28910, -28214, -25897, -23884, -19229, -15920, -13886, -8833, -3998, 
    -1387, 4836, 7708, 12720, 17260, 20691, 22162, 26310, 28549, 28171, 
    30900, 30503, 30701, 29237, 28553, 27077, 24490, 20059, 18711, 12876, 
    8660, 3528, 1780, -5478, -6683, -11280, -15205, -19578, -22929, -26382, 
    -27304, -30051, -31842, -31927, -31153, -30559, -29702, -26158, -24453, 
    -20813, -17597, -13634, -8951, -5522, -1220, 4792, 9012, 12903, 17485, 
    19032, 22125, 26314, 27405, 29775, 31310, 29929, 29808, 31020, 27060, 
    26699, 23978, 20623, 18123, 12889, 8938, 5569, 437, -2806, -6524, -11689, 
    -17002, -18414, -22319, -24720, -26203, -27636, -31292, -30787, -30835, 
    -28643, -29001, -26996, -23882, -21058, -17417, -13910, -11530, -6422, 
    -2336, 3293, 8122, 11828, 15449, 17883, 21940, 24681, 27710, 28485, 
    28961, 31002, 31110, 29857, 28023, 26882, 23044, 22018, 17837, 15044, 
    9737, 4362, 1395, -2748, -6584, -10285, -16797, -19076, -22304, -25526, 
    -26804, -28745, -31730, -31657, -29267, -29347, -28612, -26617, -26195, 
    -21659, -17166, -13300, -9394, -5751, -1238, 3638, 6842, 11711, 15269, 
    19356, 21408, 23980, 28086, 30391, 31304, 30410, 29862, 29821, 29504, 
    26292, 24000, 22729, 19112, 14708, 11863, 7220, 807, -2477, -7847, 
    -11013, -15815, -17509, -21574, -24737, -27273, -28021, -30810, -29928, 
    -32292, -31281, -29821, -26830, -24056, -22193, -18157, -14849, -11238, 
    -6415, -1013, 1372, 6162, 10269, 14704, 17902, 22402, 23131, 26371, 
    29660, 30860, 29317, 31473, 29977, 30162, 25977, 24456, 22664, 19413, 
    16785, 11656, 7436, 1705, -443, -6307, -8905, -13768, -18361, -22348, 
    -23848, -26224, -28947, -29005, -29839, -31145, -30860, -28728, -28471, 
    -25673, -21154, -18729, -15185, -9723, -7947, -4461, 1488, 5588, 10416, 
    14470, 18017, 20930, 25617, 27468, 28669, 28835, 30402, 30653, 29438, 
    30044, 26913, 24197, 22851, 19529, 16249, 10283, 7787, 2163, -1767, 
    -6507, -8831, -14359, -16575, -22045, -24857, -25783, -28834, -28560, 
    -31169, -30324, -30118, -30267, -27311, -23857, -21345, -18035, -15482, 
    -10315, -7515, -1858, 2094, 5905, 9999, 15388, 16449, 20093, 23892, 
    25445, 28467, 29144, 30514, 30947, 29987, 28976, 27029, 23804, 22723, 
    18543, 15091, 12850, 6649, 4374, -2745, -4444, -9751, -13796, -18310, 
    -20980, -23744, -27408, -29552, -29045, -29990, -31223, -29469, -29662, 
    -27964, -23882, -22138, -20371, -17387, -12018, -9205, -1987, 945, 5604, 
    8559, 13120, 16984, 21168, 24118, 25960, 28499, 29970, 30359, 30704, 
    30452, 28318, 27477, 26678, 22756, 19987, 15486, 11471, 6941, 3785, 
    -1088, -5970, -8896, -13103, -17688, -20822, -23883, -26206, -29324, 
    -29217, -31627, -29886, -30677, -31302, -27161, -27147, -21953, -20497, 
    -17476, -11898, -8509, -5340, 1453, 4592, 7774, 13809, 17513, 20032, 
    23760, 25441, 29716, 30413, 30076, 31921, 30295, 28391, 26768, 26953, 
    22699, 20009, 16331, 12558, 9036, 4961, -828, -2902, -10307, -11486, 
    -16740, -21618, -22722, -27144, -28588, -29379, -30983, -30768, -30574, 
    -29238, -26672, -26951, -23169, -18642, -17739, -12075, -10359, -3055, 
    -1190, 3559, 7522, 14199, 16065, 20618, 21751, 26719, 27475, 28842, 
    32103, 29116, 30793, 29266, 28007, 26110, 25205, 20330, 17095, 13078, 
    9002, 3938, -226, -4038, -8618, -11839, -16713, -19278, -22284, -26746, 
    -26655, -28386, -30349, -29904, -30822, -28953, -27277, -26168, -23903, 
    -20412, -17137, -11619, -8761, -3588, 573, 4767, 7298, 12439, 16354, 
    18696, 22337, 25006, 27301, 28588, 31899, 30804, 31821, 31087, 28157, 
    27697, 25306, 21269, 17292, 13266, 9995, 5052, 430, -2536, -8277, -13139, 
    -17635, -19102, -22643, -26385, -26607, -28908, -30449, -31586, -30683, 
    -28842, -29057, -26225, -21944, -19723, -17212, -14484, -9676, -5402, 
    158, 2652, 9075, 12504, 15332, 20175, 22874, 26433, 27097, 29497, 29571, 
    29922, 30115, 30019, 28194, 25747, 22781, 22066, 17396, 13309, 9802, 
    6202, 215, -4008, -6358, -11110, -14466, -20650, -23674, -24667, -27080, 
    -29597, -29757, -30560, -31910, -29357, -28281, -26313, -24999, -21063, 
    -16571, -14631, -9684, -5167, 347, 3105, 8042, 10675, 15547, 20048, 
    22535, 25298, 28028, 28741, 29329, 32097, 30645, 29253, 27244, 27687, 
    24287, 22655, 19291, 15355, 11264, 4989, 441, -2651, -6931, -12948, 
    -15127, -18627, -23400, -23931, -26202, -29365, -30134, -31624, -30536, 
    -29049, -28385, -26940, -24507, -21450, -17475, -14636, -10129, -6430, 
    -598, 3366, 8092, 12632, 15610, 19714, 22751, 25513, 27437, 30851, 30701, 
    30929, 30282, 30101, 29809, 26247, 23637, 23017, 16496, 13386, 10789, 
    6337, 3167, -2538, -6773, -9807, -14296, -17886, -20711, -25536, -27953, 
    -28291, -29336, -28907, -30534, -30803, -28109, -28163, -24349, -22006, 
    -19326, -15672, -10356, -7382, -1941, 2558, 7689, 9212, 13803, 18546, 
    21335, 24648, 26809, 30062, 30916, 31400, 32104, 30352, 29217, 27206, 
    24347, 22036, 18920, 15646, 11689, 6283, 3362, -2483, -6841, -9999, 
    -14370, -17780, -20497, -25672, -27639, -28997, -31514, -30326, -30730, 
    -31080, -29562, -28296, -23402, -20603, -20423, -15728, -11156, -6624, 
    -1734, 2011, 6629, 10037, 13128, 18593, 19716, 24697, 25666, 29100, 
    28752, 30025, 31967, 29964, 29428, 26172, 24774, 21703, 18777, 14113, 
    9784, 6388, 1990, -819, -4776, -10501, -13819, -18429, -21813, -25238, 
    -25040, -28806, -29033, -32005, -31656, -29064, -29283, -26986, -25785, 
    -22470, -20180, -14142, -10926, -7455, -4379, 1190, 6480, 10527, 14222, 
    19054, 19989, 22925, 26605, 28311, 31762, 31444, 29897, 30385, 29448, 
    27587, 26081, 23069, 20208, 15660, 11593, 8226, 3050, -681, -5402, -9740, 
    -13576, -17703, -22040, -24660, -26422, -29855, -31428, -30092, -31225, 
    -30482, -29207, -28795, -24389, -22144, -17969, -14687, -12039, -9056, 
    -3445, 944, 6648, 10943, 13613, 18071, 21468, 25542, 26276, 29886, 30005, 
    29553, 31246, 29543, 30569, 28296, 26131, 21702, 19775, 16388, 11194, 
    9328, 4287, -2143, -6434, -9238, -14150, -18459, -21540, -25039, -27557, 
    -28352, -28771, -29210, -30608, -30517, -30657, -27807, -25700, -22819, 
    -18258, -15544, -12130, -9814, -3807, 417, 3843, 9652, 13138, 17896, 
    20627, 23973, 25292, 27955, 29529, 30905, 29892, 29935, 29524, 27817, 
    26464, 22091, 21498, 16272, 13271, 8367, 4929, -684, -6057, -9875, 
    -13244, -16787, -21049, -23939, -24471, -27592, -29363, -31903, -30870, 
    -32197, -30726, -27716, -26524, -23171, -20705, -15278, -11437, -7239, 
    -5419, -680, 4665, 7571, 13345, 15972, 20307, 23120, 25998, 27389, 28984, 
    30970, 29808, 30678, 30580, 28429, 25237, 22425, 20273, 15842, 12890, 
    9837, 5158, 236, -3217, -8666, -13584, -17968, -19521, -21386, -26601, 
    -28188, -27967, -28626, -30116, -30280, -28887, -27426, -26178, -24059, 
    -20438, -17405, -12855, -8110, -5067, -314, 4682, 8256, 14183, 16939, 
    20905, 22481, 25871, 29042, 28827, 30739, 31179, 30758, 29960, 26970, 
    25165, 24138, 19820, 16252, 13687, 8838, 5087, 1440, -4214, -7664, 
    -11780, -16005, -20250, -24409, -25749, -26522, -30861, -30942, -30802, 
    -30630, -30205, -28497, -25562, -22157, -20496, -15959, -12727, -9910, 
    -4413, -590, 1960, 7766, 11296, 14942, 18884, 22066, 25968, 28142, 28363, 
    29501, 31554, 31763, 30841, 27565, 27424, 25431, 20958, 16935, 12517, 
    8387, 5203, 286, -2599, -7823, -11008, -16370, -19984, -20968, -25758, 
    -27304, -28930, -31353, -30087, -31167, -29582, -29489, -26726, -25411, 
    -19483, -16565, -13547, -10005, -4955, -1127, 2394, 7371, 11297, 14380, 
    18381, 21972, 25297, 27709, 28108, 28821, 30437, 32389, 30692, 28574, 
    25033, 24013, 21091, 18587, 14702, 11001, 6320, 6, -2294, -7209, -10850, 
    -14554, -19905, -22393, -26054, -27469, -29531, -29720, -30064, -30557, 
    -29543, -28549, -25131, -24301, -21090, -19112, -13789, -9441, -5406, 
    -680, 3115, 8288, 11557, 15154, 19018, 23451, 24418, 28197, 29760, 30171, 
    29466, 30190, 29475, 30436, 26868, 23256, 20954, 17900, 15770, 9780, 
    7107, 2975, -2324, -5546, -11232, -15914, -19599, -22737, -25071, -25815, 
    -28601, -30991, -31013, -31528, -31290, -28446, -25737, -23831, -20773, 
    -18401, -13782, -9473, -7300, -1194, 720, 5922, 10596, 14928, 18772, 
    21679, 24672, 28298, 27892, 30156, 30200, 30677, 31552, 29440, 26754, 
    26197, 21170, 17357, 15751, 12052, 6953, 3489, -3433, -7299, -11004, 
    -15189, -17343, -22753, -24201, -27297, -27950, -29820, -30957, -31081, 
    -30131, -28470, -26528, -25479, -22079, -18898, -16248, -10515, -5591, 
    -2634, 945, 5007, 10234, 14800, 16357, 21390, 24963, 25262, 28366, 30797, 
    31382, 32543, 31548, 30427, 28455, 25161, 22206, 18991, 15479, 11986, 
    6410, 3402, -1563, -5806, -10908, -13424, -16717, -21311, -22490, -26432, 
    -29728, -30658, -31542, -32553, -28891, -28500, -27778, -25174, -22364, 
    -18852, -15657, -11577, -6906, -4107, 632, 7045, 9467, 14755, 17009, 
    20915, 23910, 26383, 27398, 29875, 31575, 31885, 28877, 27917, 27394, 
    25896, 21894, 19603, 16308, 11332, 9093, 3931, -1264, -4825, -9244, 
    -14018, -18131, -20915, -23478, -26182, -29406, -29454, -30782, -29030, 
    -30419, -29634, -26284, -25374, -24250, -20203, -17215, -10196, -7483, 
    -3561, 2266, 5047, 9525, 12524, 18354, 21008, 23449, 26976, 29001, 28310, 
    31304, 31754, 30130, 29512, 26894, 26512, 22190, 21036, 15441, 12441, 
    9485, 4767, -438, -5575, -9701, -13408, -18651, -20090, -23113, -26194, 
    -26778, -30834, -29932, -29996, -28657, -29519, -29490, -26227, -24249, 
    -21431, -17484, -10611, -8524, -5718, 811, 4977, 8722, 13636, 15215, 
    21513, 22218, 26725, 28903, 29262, 30823, 29843, 29592, 30215, 26711, 
    27028, 21840, 20540, 16346, 12763, 9412, 2688, -822, -5940, -10209, 
    -13631, -16152, -19873, -23384, -27128, -27683, -28821, -31069, -32089, 
    -31266, -27857, -27355, -25036, -23263, -18721, -16567, -12999, -8712, 
    -5228, 1159, 3963, 8492, 11791, 17545, 19502, 24021, 26114, 29089, 28963, 
    29336, 30939, 32033, 29026, 26633, 24834, 24109, 20081, 17280, 12440, 
    8762, 5243, 459, -4040, -9806, -12037, -15934, -21057, -23146, -27639, 
    -28769, -28881, -31344, -31192, -30283, -28503, -26893, -25879, -23954, 
    -21179, -17192, -12926, -8865, -5320, -1847, 3020, 7257, 13499, 15409, 
    18580, 22470, 24324, 28509, 28471, 29575, 29767, 30318, 29509, 27650, 
    27158, 24587, 19606, 16838, 13667, 9335, 5084, 1388, -2269, -8181, 
    -12884, -16435, -18046, -23025, -23832, -27966, -29613, -29316, -31087, 
    -29620, -30416, -28903, -26416, -24717, -19906, -16477, -12910, -9315, 
    -5795, -1106, 3704, 7435, 11653, 15357, 18277, 24032, 24403, 26934, 
    29363, 30217, 32188, 31101, 30140, 26799, 28060, 25723, 21496, 19003, 
    13718, 10415, 6261, 2519, -4075, -7680, -12195, -14863, -18457, -23025, 
    -24723, -27695, -28273, -29864, -29302, -30282, -28793, -28493, -26576, 
    -25796, -21686, -17660, -13135, -11656, -5158, -124, 2379, 8352, 11130, 
    16113, 18486, 21973, 26299, 26353, 28957, 29487, 31241, 29525, 29740, 
    29040, 25754, 25600, 20928, 18289, 14978, 11653, 5362, 2331, -3440, 
    -6049, -10311, -15253, -18502, -22584, -25450, -26906, -28702, -30156, 
    -30627, -31636, -30292, -27760, -27974, -26174, -22927, -17016, -14274, 
    -9308, -7095, -1418, 3390, 8377, 11122, 14817, 19554, 22322, 25234, 
    28024, 28640, 30209, 31244, 30062, 30461, 27514, 25856, 25668, 21009, 
    17422, 15062, 9596, 7133, 1796, -2036, -5232, -9397, -15641, -19689, 
    -23043, -23706, -27182, -28389, -29393, -30039, -31213, -31831, -27585, 
    -26073, -24831, -22931, -18470, -14995, -11618, -8005, -1209, 2637, 6579, 
    12265, 14777, 17965, 20735, 25150, 27081, 28123, 28834, 30652, 29953, 
    30568, 28044, 26619, 24377, 20222, 19289, 15883, 11277, 8523, 2629, 
    -1637, -5099, -11408, -15162, -18766, -22829, -25021, -27700, -29314, 
    -31294, -31089, -28877, -29008, -29604, -28084, -24437, -22132, -17633, 
    -15768, -12083, -8338, -4047, 1734, 5836, 9662, 13265, 19075, 21643, 
    24432, 26092, 28915, 29239, 31585, 31306, 30357, 28434, 27050, 25883, 
    22699, 18368, 14735, 12279, 5561, 3117, -870, -5435, -10739, -13832, 
    -17621, -22858, -25180, -26468, -27921, -31501, -31739, -31492, -30843, 
    -28985, -26651, -25808, -20800, -19304, -15382, -11467, -6944, -2928, 
    309, 5752, 8755, 14101, 18210, 21935, 22568, 26751, 29535, 30776, 29463, 
    31331, 29792, 28392, 28663, 24930, 22757, 18931, 14325, 11284, 7516, 
    3171, -251, -6472, -10653, -14807, -16149, -20737, -24249, -25986, 
    -28881, -28815, -30105, -30854, -30306, -29034, -26496, -26740, -22118, 
    -18601, -15738, -12266, -7550, -2672, 1427, 4792, 9612, 14500, 18258, 
    21358, 22393, 24974, 28026, 29443, 29362, 31533, 29554, 29239, 27069, 
    26260, 21976, 19669, 16788, 12443, 7833, 5016, 82, -6017, -9136, -11534, 
    -17297, -21016, -23577, -25734, -28268, -29111, -30715, -30713, -31711, 
    -29104, -28804, -25202, -22153, -19449, -15454, -13648, -8232, -4902, 
    -967, 3884, 8207, 12795, 17580, 20768, 24099, 26897, 27851, 30232, 30785, 
    30859, 29665, 29239, 28322, 24615, 22470, 21193, 17192, 13679, 8977, 
    3659, 197, -4849, -8516, -12338, -17001, -20668, -23294, -26855, -28279, 
    -30332, -29837, -31506, -29958, -30469, -27738, -26927, -23625, -20541, 
    -17556, -12716, -8875, -3222, -107, 5640, 6957, 11785, 16898, 19894, 
    22638, 25492, 27777, 29825, 29435, 30025, 29553, 30119, 29804, 25136, 
    23569, 19422, 17950, 11982, 7933, 4104, -272, -2868, -10061, -13014, 
    -17977, -18348, -24177, -25625, -27224, -29334, -30483, -31132, -31134, 
    -29072, -28823, -26260, -22952, -19270, -16292, -14029, -7456, -4178, 
    -1595, 3383, 9197, 11903, 15972, 18519, 22130, 27261, 28743, 29921, 
    30167, 29529, 29605, 29500, 27830, 26276, 23826, 19872, 17486, 12107, 
    10385, 5026, 612, -3516, -9024, -12668, -16763, -20287, -24177, -24931, 
    -27446, -29218, -30661, -32043, -30810, -30160, -28960, -26356, -23060, 
    -20037, -17460, -14332, -10412, -5895, -498, 2719, 9306, 11637, 15609, 
    19096, 22577, 25940, 28600, 30623, 30307, 29116, 30243, 30315, 28658, 
    27557, 24512, 20365, 17826, 13420, 11343, 5280, 1576, -3139, -7717, 
    -12549, -16522, -19430, -23194, -24824, -26267, -29663, -29617, -29390, 
    -31683, -30349, -28006, -26860, -23331, -19712, -16462, -13066, -10456, 
    -6407, 280, 3762, 7594, 11393, 15319, 19170, 21641, 24324, 28010, 29183, 
    29680, 30656, 30576, 30317, 27922, 25129, 22872, 20450, 18136, 13724, 
    10285, 6048, 1863, -4148, -7625, -11467, -15056, -17838, -22520, -25257, 
    -28785, -29395, -30682, -30735, -32592, -29323, -29180, -27575, -23673, 
    -20815, -17678, -15556, -9579, -6606, -1674, 2297, 7224, 11003, 14355, 
    18883, 21765, 24509, 28097, 29912, 30446, 30798, 30384, 28602, 28425, 
    26319, 24359, 20639, 17443, 14569, 10265, 6658, 2523, -3401, -5953, 
    -11444, -14698, -18482, -22824, -23442, -26181, -29150, -30980, -29634, 
    -29639, -30376, -30248, -28756, -23217, -21825, -19306, -13385, -11446, 
    -5919, -432, 2128, 6757, 10656, 14225, 18225, 23203, 25406, 25661, 28350, 
    30625, 30657, 31682, 31629, 28329, 26734, 23270, 23082, 18872, 14403, 
    10701, 7705, 1375, -2456, -6231, -10209, -15180, -19439, -22607, -23380, 
    -26971, -29292, -29142, -30199, -31428, -31701, -28787, -28003, -25348, 
    -21605, -20112, -15780, -12331, -6236, -3523, 1675, 5812, 9402, 14884, 
    17748, 22395, 25616, 25407, 27976, 30715, 31381, 30030, 31557, 28262, 
    25778, 25659, 22054, 19730, 16785, 11326, 7837, 3067, -808, -6098, -9763, 
    -14787, -18331, -21055, -22543, -26575, -27914, -29581, -31377, -30076, 
    -29847, -27939, -27351, -25731, -22373, -18848, -15399, -11966, -6617, 
    -3652, 1446, 4420, 8980, 14305, 18738, 21515, 23874, 26406, 29237, 30139, 
    31200, 30651, 30731, 28250, 26110, 25120, 23094, 18655, 14788, 11796, 
    7845, 3337, -1286, -4983, -9857, -13909, -17217, -21352, -24305, -25940, 
    -29139, -29808, -31092, -31013, -29469, -29053, -27228, -24126, -23418, 
    -20024, -16802, -13239, -8192, -3426, 1334, 5764, 9413, 13439, 17118, 
    20058, 24828, 27529, 27796, 30957, 31691, 31018, 30712, 29965, 26797, 
    24729, 22800, 20291, 17683, 12723, 8433, 3923, -381, -4537, -9739, 
    -13280, -18265, -18947, -23657, -27337, -28603, -29571, -30945, -30812, 
    -30276, -28688, -28714, -25046, -23090, -18749, -16824, -12622, -7890, 
    -3615, 1295, 4842, 9927, 12875, 18203, 19507, 22964, 26538, 27853, 31391, 
    29962, 30154, 30523, 28797, 27646, 25448, 23117, 20059, 14930, 12364, 
    9439, 3643, -432, -3685, -8439, -12676, -17972, -19464, -22559, -24814, 
    -28540, -30782, -31612, -30461, -29970, -29716, -28459, -25304, -23231, 
    -19144, -16512, -12503, -8205, -5487, -401, 3845, 7446, 12913, 17957, 
    19786, 22960, 24540, 29702, 30502, 29781, 29687, 32201, 30676, 27217, 
    25738, 23760, 19550, 17446, 12506, 8575, 4545, -934, -3897, -9444, 
    -14000, -15472, -20150, -22454, -26213, -28132, -30162, -30722, -29707, 
    -29642, -29580, -29672, -27277, -22403, -20156, -18029, -12599, -9950, 
    -3958, 314, 3737, 8215, 13169, 16803, 21031, 24592, 26072, 26537, 28524, 
    28896, 30518, 30291, 29579, 28111, 26467, 21922, 20028, 16730, 14192, 
    9406, 5918, -28, -3280, -6389, -13191, -15486, -19039, -23097, -25178, 
    -27919, -27896, -30912, -31596, -31891, -28483, -28319, -25483, -23228, 
    -21318, -18123, -13521, -9393, -6436, -1063, 5047, 7824, 11661, 15425, 
    19044, 22672, 25066, 27971, 28632, 31138, 30959, 30035, 31144, 28187, 
    25661, 23167, 21298, 17381, 14868, 9388, 5570, -394, -2824, -8148, 
    -10112, -16234, -18758, -21873, -24137, -26921, -29026, -30880, -31946, 
    -29667, -30284, -28960, -26671, -24665, -21217, -17661, -13066, -11411, 
    -5557, -1390, 4315, 7695, 11214, 15961, 17761, 24020, 25351, 26694, 
    28521, 30829, 32150, 30069, 31147, 28781, 26340, 24616, 20082, 18588, 
    12839, 10766, 6470, -54, -3406, -6064, -11133, -15300, -19163, -23319, 
    -24769, -28045, -29769, -30544, -30695, -30628, -28326, -29970, -27620, 
    -24476, -22280, -18021, -14628, -10113, -4855, -1321, 3631, 7733, 11764, 
    14901, 19865, 23121, 25661, 26869, 28973, 29731, 29389, 31850, 30381, 
    28816, 26406, 24865, 21510, 18447, 13165, 9584, 7349, 2719, -3287, -5828, 
    -10855, -16001, -20192, -21918, -24756, -26453, -29583, -28893, -30118, 
    -31432, -30632, -28697, -26503, -24131, -22428, -17983, -14743, -10740, 
    -6049, -1731, 2214, 6292, 11873, 12997, 18826, 21999, 23592, 25364, 
    28362, 30223, 30195, 31123, 31579, 28169, 25502, 23700, 20976, 17826, 
    13659, 11452, 6420, 2070, -1923, -7361, -9259, -14796, -17390, -20362, 
    -24764, -27601, -30120, -30105, -29656, -29440, -29214, -29024, -26928, 
    -24488, -20841, -18883, -14432, -11254, -6541, -2539, 3051, 5467, 9801, 
    14989, 17698, 22397, 24916, 27520, 28305, 29881, 31044, 30245, 30025, 
    28592, 27539, 25195, 22439, 17863, 15649, 11794, 6553, 3954, -2314, 
    -4618, -11901, -12505, -17408, -21106, -24227, -26859, -28844, -28776, 
    -30940, -31026, -30127, -28064, -26931, -25836, -22252, -20510, -15474, 
    -11605, -7114, -3956, 1542, 6198, 9880, 13265, 16307, 21363, 23248, 
    27397, 29125, 31170, 30578, 30622, 30860, 28327, 27146, 26753, 23188, 
    18968, 16755, 10644, 6367, 4219, -2191, -5305, -11099, -12419, -17014, 
    -20327, -25407, -26581, -28661, -28672, -31636, -31206, -29578, -28593, 
    -27890, -26474, -22294, -19478, -15230, -11853, -8456, -4361, 896, 4813, 
    8995, 13827, 17418, 19948, 23930, 26462, 28719, 29243, 30647, 30470, 
    30957, 29826, 26768, 25126, 21447, 19308, 16812, 11373, 8317, 3141, 
    -1221, -6392, -10420, -13050, -17607, -19880, -24329, -26418, -28611, 
    -28928, -31453, -30705, -31346, -30589, -28383, -25686, -22478, -19690, 
    -17508, -12675, -8168, -4477, 1748, 4653, 9775, 13157, 16827, 21697, 
    22728, 26482, 28691, 30367, 31039, 29880, 29425, 29513, 27983, 25836, 
    23507, 18658, 17446, 13124, 8818, 3920, -928, -5095, -8797, -13040, 
    -16876, -20299, -23577, -25807, -28659, -30162, -28895, -30152, -29706, 
    -29100, -28233, -25232, -24307, -21958, -16683, -12509, -7971, -4232, 
    -910, 3873, 9980, 13470, 18277, 19009, 22915, 25838, 28374, 29028, 31509, 
    29545, 29887, 28413, 28193, 24927, 25086, 19804, 15355, 12454, 9239, 
    4861, 703, -4501, -8478, -12656, -16494, -20115, -22262, -24975, -27187, 
    -29431, -32133, -30635, -29743, -30067, -29155, -25518, -23834, -19906, 
    -17312, -12950, -9752, -4059, 62, 4145, 6952, 12242, 16764, 19809, 22711, 
    25075, 28054, 29272, 31353, 30968, 30583, 30667, 28460, 27123, 23306, 
    19761, 16477, 14227, 8949, 4677, 606, -2195, -7899, -11903, -16705, 
    -19537, -23963, -26449, -26745, -31189, -29521, -30812, -31261, -29729, 
    -28140, -26112, -22289, -19702, -17278, -14892, -10137, -4665, 483, 3321, 
    9343, 12589, 14395, 19319, 21681, 24172, 27830, 28634, 30470, 32280, 
    31501, 29865, 27263, 26595, 24315, 21862, 16626, 12867, 9515, 7293, 858, 
    -4651, -8662, -12992, -17214, -20751, -21829, -25379, -26686, -29614, 
    -30581, -30361, -30641, -29491, -28781, -26779, -23565, -21388, -18667, 
    -15186, -9166, -5392, -261, 3169, 5626, 11816, 16348, 19938, 22744, 
    25177, 25993, 30708, 29914, 29415, 29349, 29906, 27397, 26113, 25130, 
    22122, 18575, 13927, 10651, 6741, 1015, -3216, -7432, -11643, -16631, 
    -18969, -21093, -25632, -26015, -30273, -31678, -31981, -30967, -29886, 
    -27840, -27028, -22492, -20155, -17721, -13479, -11669, -4993, -2308, 
    1060, 5940, 10846, 16606, 17597, 22063, 24624, 26630, 30047, 30034, 
    30392, 31465, 28422, 28735, 26554, 26104, 20359, 17555, 14365, 11498, 
    6558, 1579, -3064, -5826, -10244, -14331, -17300, -21277, -25240, -26704, 
    -29513, -30752, -32190, -31267, -30868, -29513, -26158, -24666, -21676, 
    -18603, -15669, -9705, -6769, -3040, 612, 5733, 11496, 14312, 18701, 
    21733, 22973, 25370, 29614, 30061, 30250, 32353, 28888, 28324, 27571, 
    23473, 23065, 19308, 13432, 9510, 7584, 3097, -2117, -5239, -10130, 
    -14760, -18774, -20223, -23750, -27793, -29324, -28957, -30128, -31777, 
    -30651, -29060, -27691, -24038, -22970, -18516, -14509, -10172, -6717, 
    -3102, 481, 7214, 9391, 14088, 17758, 22582, 23823, 27682, 28585, 31097, 
    30198, 30500, 28911, 29677, 25868, 24741, 22469, 18791, 15307, 10458, 
    6951, 2849, -1522, -6036, -10167, -14714, -18858, -20597, -24206, -25791, 
    -29379, -30809, -29057, -29982, -30838, -29995, -26760, -25669, -22895, 
    -18547, -15404, -12388, -7424, -3145, 2067, 5341, 9708, 14209, 19170, 
    22300, 24881, 27805, 29103, 30847, 31001, 31136, 29419, 28286, 26558, 
    26637, 21756, 19192, 15676, 10796, 6288, 2690, -1091, -5283, -9712, 
    -14453, -17893, -21298, -23963, -27242, -27309, -29314, -30568, -30734, 
    -28466, -28696, -27184, -26212, -21458, -19475, -16056, -11421, -9125, 
    -4984, 1232, 6359, 9394, 13716, 17782, 20865, 24001, 26084, 28947, 29528, 
    31722, 30995, 29751, 27723, 28788, 25653, 22876, 21320, 17002, 12547, 
    7803, 4751, -1050, -4703, -10118, -13728, -16523, -21031, -23483, -26775, 
    -27263, -30410, -31241, -29670, -29897, -30609, -27895, -25998, -23510, 
    -19976, -17680, -11599, -9012, -3499, -1068, 5036, 8057, 11296, 15816, 
    21578, 22764, 24425, 27320, 31403, 29931, 29825, 30045, 30006, 26422, 
    26121, 21634, 20282, 16085, 12450, 9849, 4712, -371, -3543, -8945, 
    -14138, -17436, -20414, -22000, -26479, -27548, -29332, -31423, -30134, 
    -32148, -30007, -27364, -26027, -23483, -21178, -17272, -13335, -8814, 
    -4283, -286, 4180, 8644, 13346, 16039, 19973, 23775, 25155, 28201, 30273, 
    29176, 31660, 31198, 29345, 27676, 26455, 23692, 21102, 16405, 11990, 
    9806, 4035, 495, -3603, -8276, -12247, -15941, -18753, -23404, -26578, 
    -28227, -28278, -30906, -29498, -31928, -31048, -28496, -25480, -23659, 
    -21966, -15924, -14017, -7320, -4879, 5, 2570, 7930, 12454, 16372, 19444, 
    21622, 25514, 27663, 29486, 30442, 30089, 30432, 28756, 27619, 26266, 
    23126, 20830, 16663, 13350, 10344, 6140, 322, -3083, -7942, -12636, 
    -16294, -19053, -21218, -26339, -27505, -29273, -30916, -29285, -31284, 
    -30453, -28481, -25515, -23769, -20600, -17888, -13267, -8917, -3676, 
    -746, 3760, 7872, 10053, 15663, 19163, 22511, 25258, 27928, 28401, 30889, 
    29945, 30011, 28944, 26827, 27163, 23291, 21234, 18265, 14870, 9665, 
    4346, 1167, -2591, -8993, -12272, -15452, -19943, -22941, -23495, -28334, 
    -29491, -30754, -30247, -30098, -29825, -28557, -27744, -24678, -22665, 
    -18480, -14827, -9299, -5431, -1090, 3065, 7086, 11403, 15113, 19023, 
    22597, 24069, 27595, 27804, 29881, 31604, 31845, 30337, 28196, 25299, 
    24130, 21599, 16771, 13793, 10688, 4284, 326, -3844, -7889, -10634, 
    -14557, -19706, -22403, -25853, -26077, -28705, -30767, -29837, -30756, 
    -30942, -28702, -27353, -22848, -22283, -17733, -15289, -10838, -5881, 
    -1032, 3157, 5400, 10359, 15309, 18255, 22756, 24294, 26947, 29021, 
    30635, 30311, 31602, 30724, 29342, 26764, 24563, 20753, 18127, 14359, 
    10308, 6978, 1216, -3033, -6762, -10619, -15316, -18906, -23118, -24478, 
    -27743, -29451, -29948, -29934, -31640, -31568, -28662, -28079, -24716, 
    -20744, -18975, -14720, -11182, -6005, -2068, 2010, 5993, 10577, 14718, 
    19391, 21502, 25442, 26917, 28650, 29744, 30612, 29861, 30189, 28167, 
    27482, 24389, 20528, 19432, 15977, 9561, 6977, 2391, -2168, -6661, 
    -12136, -13021, -17610, -21336, -23744, -27004, -27966, -31827, -29462, 
    -30806, -29496, -29447, -26603, -24629, -22303, -18196, -16097, -11833, 
    -7331, -1890, 1726, 5404, 11267, 15480, 18134, 21006, 24009, 27611, 
    28342, 31444, 29163, 31070, 29739, 29842, 25682, 25686, 22926, 20301, 
    16463, 11639, 7484, 3585, -1466, -5162, -10097, -15284, -17037, -20668, 
    -25226, -26355, -28936, -31388, -31121, -32111, -30980, -29495, -28489, 
    -24089, -22683, -19145, -15512, -11609, -7732, -3179, 1301, 4400, 9938, 
    15093, 18009, 22925, 24494, 26295, 28579, 30339, 32068, 30408, 31369, 
    30003, 26109, 25975, 22916, 20161, 16724, 11626, 7807, 3465, -12, -4187, 
    -8426, -12699, -17764, -19973, -23741, -26710, -27675, -29696, -31103, 
    -30434, -30495, -29079, -27718, -26198, -21394, -19789, -16191, -10351, 
    -7423, -3435, 611, 4791, 10480, 13178, 17330, 19855, 22710, 26598, 29700, 
    30536, 30890, 29256, 29880, 30498, 28187, 26434, 24046, 20862, 17197, 
    11041, 7808, 2750, -780, -4711, -9300, -12165, -18441, -21184, -25243, 
    -25258, -27795, -29572, -30688, -32379, -29850, -29401, -27492, -24788, 
    -22859, -18648, -15781, -11143, -9606, -4768, 1933, 5727, 9410, 13862, 
    17037, 21271, 23586, 25821, 28600, 29327, 30679, 30810, 29481, 29385, 
    27309, 26007, 24436, 21057, 17675, 12450, 9919, 4892, 1349, -3886, -8687, 
    -12397, -16937, -22064, -24394, -27425, -28246, -29794, -30814, -30803, 
    -30583, -30190, -26567, -25102, -22510, -21668, -17447, -13317, -9958, 
    -4669, -660, 3413, 8812, 12114, 16405, 20701, 23526, 27040, 26553, 29530, 
    30847, 31268, 30738, 29865, 29268, 26727, 23654, 19793, 16659, 13577, 
    9014, 4614, -23, -4327, -9895, -12956, -15841, -19170, -23452, -26251, 
    -28343, -29544, -31029, -30379, -30729, -29752, -29361, -26111, -24427, 
    -22333, -18150, -13722, -7970, -4849, -1317, 3945, 9368, 12676, 16043, 
    18743, 23337, 25472, 26887, 29973, 30835, 29999, 30661, 29315, 27219, 
    24902, 23273, 21569, 17997, 12610, 9012, 5118, -125, -4424, -8410, 
    -14054, -14860, -21016, -22464, -26990, -29402, -29384, -30882, -30872, 
    -29842, -31335, -27434, -26638, -24514, -21146, -16804, -14276, -9056, 
    -4931, 189, 2600, 8741, 11524, 16491, 18412, 23232, 25414, 28234, 29091, 
    31399, 31433, 30053, 29194, 28748, 27121, 25013, 21474, 17588, 14964, 
    7873, 3695, 2214, -4724, -6421, -11020, -17302, -20903, -21623, -25518, 
    -27106, -28914, -29831, -30346, -30624, -30548, -30015, -26120, -23294, 
    -22275, -17143, -14517, -11604, -6401, -1947, 3489, 7230, 11876, 16380, 
    19991, 21175, 23686, 27049, 29983, 31540, 30930, 30685, 28926, 28000, 
    26868, 24494, 20925, 18774, 14280, 9366, 6021, 1025, -3103, -8350, 
    -12545, -15667, -18835, -22164, -24188, -27740, -28733, -31562, -30791, 
    -31311, -30449, -28937, -25881, -25584, -22918, -19368, -14280, -10056, 
    -5362, -2981, 3703, 7126, 10540, 15888, 19290, 22453, 23681, 27398, 
    27482, 30746, 31255, 30017, 30965, 27865, 25393, 23943, 21561, 18069, 
    15697, 9015, 6917, 497, -2105, -7184, -10874, -14651, -18654, -21920, 
    -24811, -25985, -29039, -31260, -30650, -30218, -29952, -28211, -26982, 
    -25123, -22559, -18132, -14991, -10134, -5207, -643, 2261, 5728, 10976, 
    15847, 17063, 21525, 23651, 26942, 29750, 30790, 31360, 29052, 29805, 
    28630, 26782, 24993, 20565, 19585, 15893, 12678, 7554, 2682, -1214, 
    -6259, -10735, -13819, -17871, -21064, -24098, -25983, -28697, -28664, 
    -31411, -30771, -30173, -27421, -26628, -26598, -21090, -18505, -13625, 
    -11527, -6469, -2860, 2748, 7338, 10631, 14431, 18247, 20315, 23952, 
    27711, 28818, 29232, 30212, 31931, 31617, 29760, 28699, 24853, 21078, 
    17845, 15674, 9864, 8841, 4408, -1270, -6555, -10215, -14089, -17437, 
    -20593, -23183, -25954, -28695, -29925, -31103, -31456, -29627, -28941, 
    -26710, -25412, -23223, -19360, -14650, -12416, -6862, -2875, -111, 5599, 
    11089, 13047, 17086, 20764, 24084, 26937, 27028, 29947, 30168, 29481, 
    30644, 29251, 28165, 23690, 22675, 19003, 16514, 12709, 8233, 3424, 
    -1602, -6127, -9285, -14985, -16440, -21265, -24008, -26631, -28291, 
    -30536, -31864, -29882, -29607, -30079, -27303, -24839, -22014, -18670, 
    -17205, -12567, -7650, -3476, 649, 4216, 8309, 13989, 18718, 20770, 
    23135, 26857, 28005, 29837, 30104, 30870, 29797, 30253, 28796, 25671, 
    23017, 20754, 14699, 12785, 7692, 4068, 412, -3924, -9140, -14319, 
    -17014, -21101, -22341, -24617, -27494, -29821, -30522, -31208, -30358, 
    -29332, -26456, -26494, -21747, -19231, -16366, -13006, -8815, -4787, 
    145, 4155, 9588, 11771, 17496, 21305, 23608, 26520, 29064, 30333, 29767, 
    30660, 29675, 29737, 28128, 25908, 22910, 20909, 16323, 13264, 9517, 
    3003, -412, -4084, -10041, -12245, -18062, -19195, -24575, -25676, 
    -28081, -30382, -31018, -31789, -29648, -29206, -28262, -27090, -24371, 
    -19380, -16530, -12305, -8640, -4161, -198, 3971, 9215, 13113, 17599, 
    19462, 23140, 26728, 28715, 28950, 29714, 29763, 30725, 29981, 27780, 
    26106, 23103, 21607, 16851, 13914, 9736, 5582, -117, -3218, -7728, 
    -11901, -15306, -20010, -22267, -25458, -27326, -30249, -30129, -32461, 
    -31574, -29837, -28076, -25404, -24204, -19706, -18132, -13062, -7625, 
    -4396, -209, 3523, 8358, 11766, 16234, 20420, 21231, 26710, 27817, 29828, 
    30782, 30653, 30982, 30155, 27568, 26358, 22534, 21368, 17099, 13129, 
    8513, 6720, -203, -3463, -7785, -12796, -17363, -18731, -23523, -25705, 
    -27763, -29108, -30871, -30936, -30565, -28908, -27395, -25849, -24504, 
    -22496, -16445, -13316, -9028, -4889, -1270, 3310, 7234, 13351, 15464, 
    19786, 21652, 26142, 28329, 28496, 31133, 32107, 31151, 29058, 28868, 
    26203, 23882, 20281, 19306, 13352, 8386, 4340, 556, -2684, -7488, -12417, 
    -15672, -20129, -22676, -23726, -27997, -29212, -31127, -30227, -30862, 
    -29847, -27814, -26982, -23407, -21936, -16467, -14021, -10163, -4974, 
    -1246, 3359, 6521, 11158, 16122, 18498, 22664, 24731, 27669, 29195, 
    30576, 31228, 29443, 29328, 27770, 27128, 23073, 22730, 16881, 14338, 
    10121, 6483, 2207, -4602, -7240, -12229, -15144, -19053, -22924, -25691, 
    -27615, -28980, -30245, -30064, -31507, -31035, -27439, -27984, -23715, 
    -22022, -19105, -13356, -11668, -5790, -1588, 3513, 6353, 11961, 15080, 
    17799, 20383, 25214, 28142, 28675, 30523, 30795, 31489, 31448, 27164, 
    26814, 25501, 22195, 18655, 15664, 9957, 4916, 3064, -2196, -6995, 
    -10556, -14774, -18342, -20590, -25407, -26738, -28754, -30315, -30480, 
    -29302, -29159, -29429, -27852, -23687, -21890, -19523, -15172, -9791, 
    -6795, -3245, 1343, 6739, 10831, 15640, 17599, 21370, 26145, 26454, 
    28667, 29571, 30607, 30637, 31139, 28945, 28442, 24865, 22441, 18225, 
    14866, 10039, 8487, 2600, -2409, -5080, -11499, -14004, -18041, -20945, 
    -24411, -26075, -29270, -30123, -30007, -30028, -30779, -29648, -27034, 
    -25840, -23049, -17647, -14580, -10515, -6673, -1122, 1204, 5601, 10169, 
    14147, 18269, 19737, 23904, 28003, 28426, 30258, 29980, 30473, 29897, 
    29573, 28144, 24241, 21324, 17224, 14801, 12762, 7967, 1868, -808, -5287, 
    -9064, -13740, -16801, -21509, -25342, -27439, -28656, -31280, -30248, 
    -29053, -29430, -28145, -27585, -24853, -21519, -19398, -15114, -11146, 
    -6646, -2341, 1433, 5990, 11025, 15225, 18034, 20434, 23966, 25685, 
    28445, 29791, 31711, 29977, 29473, 28782, 27211, 23655, 23257, 18972, 
    14972, 12727, 6502, 3467, -1425, -5011, -8701, -13968, -17619, -21071, 
    -23836, -27016, -29654, -29278, -31152, -31306, -29820, -29420, -27997, 
    -25092, -23790, -19037, -17247, -11530, -8475, -2244, 2448, 5369, 9778, 
    15480, 17669, 21226, 22497, 26824, 27868, 31650, 30008, 31478, 29759, 
    30021, 28298, 24659, 22040, 19668, 15981, 11498, 8756, 5179, -2109, 
    -5263, -8536, -13799, -18545, -21439, -24249, -24615, -27881, -28351, 
    -30726, -30908, -29801, -29613, -26278, -25601, -22454, -18857, -17096, 
    -12159, -9012, -3628, 745, 3821, 9875, 11940, 16929, 19442, 24415, 25189, 
    29175, 29522, 30979, 30663, 30082, 30696, 27228, 26628, 24010, 18563, 
    17662, 12470, 7625, 4773, -1735, -3667, -8272, -13946, -17446, -21902, 
    -22814, -25674, -27781, -29619, -31008, -32114, -29992, -29419, -27409, 
    -25010, -22855, -20258, -17279, -12754, -8893, -5365, -89, 5945, 7810, 
    13913, 18263, 20195, 22086, 26935, 28784, 29591, 31799, 31341, 30015, 
    29394, 29594, 26482, 24070, 19851, 16724, 13276, 9323, 4344, -135, -3490, 
    -8879, -11908, -17296, -20002, -24333, -26239, -27983, -29439, -30962, 
    -31872, -30305, -29994, -27958, -26915, -23571, -21120, -16881, -13293, 
    -10022, -5136, -238, 2844, 7786, 11617, 16461, 18849, 22126, 25546, 
    26603, 29613, 30521, 30582, 29689, 28777, 27999, 25684, 23980, 20477, 
    17522, 13287, 9435, 6379, 1511, -3732, -8863, -11246, -16365, -20566, 
    -24362, -25640, -26561, -29879, -31495, -30060, -28911, -29370, -28399, 
    -26323, -24604, -21430, -17443, -13549, -9670, -6502, -1394, 4126, 6718, 
    12310, 14988, 19912, 23123, 24858, 27326, 28588, 29548, 30568, 29623, 
    30169, 27388, 25091, 22965, 20777, 17066, 12835, 9236, 5441, 1699, -3303, 
    -6875, -9975, -14470, -19964, -22983, -26051, -28735, -28340, -31255, 
    -30514, -29435, -29060, -28420, -27684, -24385, -19677, -17794, -15106, 
    -10595, -7060, -1082, 3383, 7919, 11845, 16594, 18531, 22027, 24688, 
    27621, 28158, 28896, 30547, 30084, 29643, 29108, 27087, 25319, 21041, 
    18703, 13885, 10208, 6597, 1119, -3735, -6729, -10807, -15809, -19992, 
    -21575, -24765, -27845, -29005, -30684, -30861, -31166, -29468, -28549, 
    -26460, -23107, -21427, -17132, -14094, -10280, -6501, -3050, 1459, 7091, 
    10399, 15376, 18433, 22011, 25397, 26175, 29657, 30657, 31870, 31872, 
    29140, 29996, 27538, 24204, 21455, 18099, 14414, 11910, 6418, 783, -735, 
    -7366, -10502, -14798, -18954, -22002, -24445, -27632, -29525, -30726, 
    -30350, -29479, -29721, -28367, -26177, -24579, -23057, -18586, -13884, 
    -12040, -7383, -2838, 2022, 6964, 10247, 15548, 18260, 22331, 26155, 
    27411, 28723, 31296, 30917, 30830, 29617, 28777, 26666, 25778, 21588, 
    17902, 15895, 9392, 6545, 1617, -3408, -6910, -11101, -13484, -16774, 
    -22408, -24413, -28063, -29566, -30085, -30373, -32266, -29878, -29121, 
    -26824, -24984, -23241, -19672, -14917, -11329, -8619, -1087, 2795, 6205, 
    9152, 14772, 18826, 23260, 24637, 27238, 28849, 30952, 30941, 31264, 
    31501, 30025, 27791, 26184, 21293, 20513, 14744, 11489, 7322, 1629, 
    -1512, -7212, -10249, -14183, -18718, -21279, -24107, -27197, -30140, 
    -28781, -31603, -30225, -31714, -29018, -27312, -25442, -21292, -18773, 
    -14757, -9758, -7223, -1740, -138, 5325, 8830, 14179, 18199, 20834, 
    24037, 27444, 29197, 30610, 30130, 29753, 30747, 30155, 27815, 26946, 
    23109, 18461, 16611, 11986, 8714, 2288, -1228, -7202, -9495, -14543, 
    -18167, -21974, -25067, -25497, -29496, -28332, -31598, -31767, -30257, 
    -28744, -28442, -25602, -21819, -20166, -16398, -12118, -6373, -4936, 
    -711, 4329, 9315, 12375, 16042, 20521, 24028, 26315, 29409, 30709, 30539, 
    31494, 29969, 30127, 28586, 24586, 22502, 19248, 17140, 10829, 6877, 
    4718, -1134, -6471, -7542, -12815, -18792, -20261, -23689, -24761, 
    -27320, -30450, -30699, -32336, -29151, -29686, -28576, -25518, -22380, 
    -20097, -17610, -12187, -8409, -4259, 1055, 5693, 8661, 12573, 17441, 
    21261, 22896, 26232, 28101, 29287, 29070, 29253, 29645, 28229, 26411, 
    25039, 22859, 19191, 15289, 13478, 9653, 3460, -1737, -3486, -9520, 
    -13609, -16352, -19553, -23910, -25638, -27432, -28468, -30591, -30843, 
    -31214, -28759, -29521, -26063, -23014, -20556, -16341, -12115, -8321, 
    -5847, -31, 3280, 8015, 11716, 16833, 20409, 23098, 25242, 26710, 29324, 
    31260, 30396, 30509, 29878, 28297, 26476, 24776, 21476, 16435, 12263, 
    8821, 3066, 63, -4024, -7602, -12747, -16013, -19407, -23153, -25591, 
    -27403, -30350, -31457, -31057, -29497, -29246, -29263, -25933, -24574, 
    -20207, -16593, -15044, -9098, -5249, -288, 3788, 8396, 12483, 16432, 
    20125, 22697, 25649, 27009, 28153, 31566, 30975, 31561, 29719, 26864, 
    24973, 22598, 20687, 17520, 13928, 8249, 5062, 505, -2863, -8734, -11778, 
    -15132, -20060, -24050, -25152, -28065, -29689, -31522, -31802, -29932, 
    -30781, -28848, -26913, -23677, -21365, -17276, -14345, -10359, -5554, 
    -811, 3013, 7015, 11431, 14984, 19668, 21888, 24599, 26221, 29669, 30077, 
    30133, 31468, 30153, 27277, 25520, 23816, 21826, 16956, 14192, 10711, 
    6068, 1286, -2913, -6514, -11574, -15699, -17747, -21349, -24909, -27964, 
    -27756, -29048, -31262, -29743, -29512, -28027, -27976, -23677, -19947, 
    -17132, -12504, -11069, -6886, -2161, 4401, 8654, 11975, 15523, 18882, 
    23185, 25590, 27158, 28856, 29319, 30436, 29508, 30258, 28984, 27260, 
    23266, 21927, 18232, 14584, 10089, 5168, 1992, -1776, -7951, -12257, 
    -15874, -19929, -22384, -24982, -26095, -28797, -30643, -31761, -29402, 
    -28459, -29204, -27634, -22815, -21207, -18175, -15195, -10795, -6071, 
    -1513, 2107, 7381, 11572, 15106, 17301, 21426, 24201, 26525, 30818, 
    28606, 29915, 29875, 29730, 30271, 27730, 25434, 22284, 17469, 15474, 
    10252, 6907, 1757, -2103, -8246, -11667, -15619, -18245, -21356, -24902, 
    -27032, -30001, -28945, -31429, -29522, -30890, -28242, -26778, -24213, 
    -20933, -17953, -14213, -11464, -6528, -3858, 505, 6684, 11758, 15456, 
    18588, 22428, 24455, 27983, 30446, 29600, 31143, 29999, 30425, 28479, 
    28484, 25461, 22696, 17720, 14455, 10460, 8243, 2375, -1089, -4928, 
    -10144, -15053, -18320, -22707, -24057, -27140, -27494, -29406, -29945, 
    -30165, -30286, -29090, -26173, -25000, -22142, -19813, -13633, -11803, 
    -7261, -2631, 2137, 6060, 10214, 13697, 17020, 20343, 23583, 27547, 
    28526, 29696, 30372, 29705, 29643, 29413, 26699, 24648, 22991, 17493, 
    15893, 11611, 8338, 3151, -1799, -4709, -11910, -15213, -19527, -20274, 
    -24509, -26509, -28660, -28944, -30918, -30645, -29934, -29735, -26375, 
    -25339, -21164, -18360, -15638, -12017, -7884, -3553, 952, 4609, 9822, 
    13955, 16494, 21185, 25464, 25664, 27932, 30477, 31462, 30219, 30392, 
    29094, 27620, 26037, 22143, 20191, 14715, 10381, 6208, 3042, -1691, 
    -5538, -9446, -15440, -18551, -21626, -24617, -25860, -28002, -30091, 
    -31083, -31765, -29980, -28079, -28157, -26284, -23348, -20396, -16563, 
    -13099, -8303, -2331, 2337, 6100, 7820, 13231, 17995, 21169, 24426, 
    25241, 29321, 30143, 30158, 30704, 29810, 29978, 27396, 25616, 22708, 
    17781, 14716, 12292, 7604, 2312, -1032, -4435, -9165, -13172, -17341, 
    -20407, -24779, -25842, -28221, -30340, -29494, -30759, -30517, -28301, 
    -27561, -26189, -22335, -21647, -17022, -10797, -8878, -5600, -148, 6037, 
    9712, 13990, 18195, 21465, 23539, 25272, 28307, 31005, 30933, 32113, 
    30415, 29498, 26517, 26364, 23136, 20639, 15271, 13201, 10021, 3701, 
    -2093, -5787, -8986, -13956, -15968, -21670, -23962, -26852, -26756, 
    -31431, -29368, -32266, -29313, -30216, -26997, -27305, -24527, -20895, 
    -16963, -13406, -9138, -3744, 85, 5472, 9676, 12927, 17306, 19180, 23275, 
    25656, 27671, 30909, 30307, 30823, 29492, 29489, 29162, 26556, 23191, 
    20810, 16998, 13347, 8598, 5332, 878, -4881, -9438, -12783, -15732, 
    -19057, -24483, -25425, -28114, -29672, -30731, -32592, -31700, -28828, 
    -29345, -25388, -23497, -21000, -17068, -13380, -8918, -4488, -1552, 
    2938, 7399, 12602, 16734, 19212, 23283, 25701, 27719, 29777, 28816, 
    29273, 31318, 29593, 28452, 25045, 23046, 20886, 17214, 13421, 9331, 
    4803, 133, -4946, -7744, -12842, -14937, -21104, -23678, -26676, -27511, 
    -30076, -29364, -31653, -31795, -29926, -28640, -26983, -23479, -20681, 
    -16713, -13857, -8042, -4747, -850, 3384, 6938, 13115, 16233, 20357, 
    23679, 26006, 27833, 29801, 30853, 30580, 29742, 29869, 28147, 26087, 
    23853, 19611, 16579, 14032, 8730, 4725, 947, -1657, -7962, -11718, 
    -14899, -19695, -21590, -24175, -26100, -29892, -29851, -31811, -31123, 
    -29248, -28466, -26399, -24471, -20395, -18281, -14870, -10374, -5740, 
    -2188, 3333, 7322, 11104, 16417, 18418, 21969, 25995, 27500, 29307, 
    30409, 30725, 31100, 31008, 28883, 26169, 23936, 22290, 17464, 14685, 
    9923, 6109, 1070, -1161, -8262, -11399, -14763, -19258, -23328, -25022, 
    -27258, -29815, -29957, -29405, -30529, -30967, -29727, -25915, -23381, 
    -20928, -18335, -13618, -10869, -5262, -3419, 2710, 8218, 11844, 14936, 
    18556, 21135, 24850, 26879, 29768, 31305, 31614, 29993, 30145, 27506, 
    27577, 24196, 21559, 17956, 16172, 11083, 5175, 2697, -3593, -6206, 
    -11273, -16535, -17873, -22478, -24867, -27513, -28218, -30747, -30123, 
    -32288, -29784, -30575, -27316, -23414, -22455, -16769, -14968, -10309, 
    -7928, -2584, 2635, 7325, 9747, 13856, 17991, 21697, 23883, 26875, 28712, 
    30034, 30351, 31236, 31750, 29551, 26194, 25286, 20402, 18981, 14692, 
    10848, 7146, 2582, -2645, -6438, -9391, -15036, -17991, -21905, -24233, 
    -27406, -29437, -31657, -29831, -31043, -28446, -30703, -27831, -24535, 
    -22172, -18686, -15228, -11110, -6766, -1247, 758, 7024, 9243, 12921, 
    17378, 21059, 24548, 26801, 29638, 31130, 29391, 30491, 28878, 30111, 
    26038, 26227, 23616, 19270, 14934, 11298, 8472, 3054, -1153, -7496, 
    -10048, -13626, -18233, -22030, -25888, -27278, -29258, -29932, -30920, 
    -30487, -30518, -28356, -28158, -26054, -22113, -19245, -15539, -11648, 
    -6082, -2467, 1635, 6909, 10131, 14007, 18083, 22089, 24036, 27346, 
    28119, 29028, 30672, 31347, 30576, 29238, 28040, 24474, 22940, 19579, 
    15433, 10761, 7714, 3096, -1914, -4646, -10453, -13190, -17316, -21233, 
    -22989, -25507, -30013, -30269, -29935, -31379, -29721, -29488, -27447, 
    -25826, -21898, -20121, -16348, -12748, -7920, -5375, 1417, 5576, 9973, 
    13423, 17044, 21784, 23956, 27265, 28518, 28302, 31182, 30832, 30493, 
    29325, 28052, 25238, 22522, 18622, 14866, 11650, 8170, 2556, -932, -4871, 
    -9295, -13282, -16530, -20634, -24628, -26917, -28973, -29672, -29066, 
    -29781, -28948, -28255, -28425, -25766, -23647, -19215, -16237, -11044, 
    -6748, -4145, 1131, 3841, 9876, 13167, 18621, 20802, 23015, 27337, 29129, 
    30386, 31681, 29677, 29427, 30096, 27971, 25028, 23075, 20195, 15873, 
    12287, 8360, 3919, -573, -5419, -7985, -11806, -16863, -19649, -23582, 
    -24498, -28587, -30017, -30583, -31306, -30582, -28793, -29428, -24232, 
    -23760, -20300, -15109, -14212, -9916, -4895, 103, 3622, 10079, 14182, 
    16821, 20881, 22802, 24122, 28200, 29505, 29341, 30459, 32136, 28915, 
    26969, 25834, 23054, 20390, 16768, 11832, 9505, 5828, 89, -3926, -8536, 
    -10999, -16627, -19801, -22825, -26288, -27793, -27772, -29849, -30878, 
    -29243, -28630, -28578, -24465, -22680, -19826, -17907, -13930, -8067, 
    -4261, -1442, 2409, 6987, 13056, 15909, 19812, 23356, 24624, 27534, 
    29530, 29385, 31359, 30021, 30347, 29682, 25464, 23223, 21491, 16339, 
    14732, 8930, 3888, 884, -3196, -8002, -12278, -15382, -19297, -21731, 
    -24446, -27400, -29461, -32131, -29912, -32263, -29776, -28443, -25998, 
    -23489, -21416, -17383, -13730, -10156, -5335, -220, 2821, 7216, 11796, 
    17468, 19525, 22172, 25456, 27829, 29232, 30938, 31088, 31956, 28000, 
    26742, 26876, 22966, 20175, 18184, 15260, 10451, 4586, 1439, -2873, 
    -7036, -11532, -14473, -19754, -22194, -25048, -28194, -28761, -31006, 
    -30639, -30074, -28954, -29530, -26293, -25140, -21705, -18212, -14604, 
    -10951, -6905, 98, 2242, 6173, 11594, 16727, 20094, 22391, 24600, 27413, 
    30361, 31843, 31402, 30457, 30608, 29237, 27540, 23885, 20439, 17061, 
    14576, 9045, 5691, 1637, -1305, -7263, -10465, -16101, -19807, -21628, 
    -25926, -25634, -30715, -30051, -30936, -31242, -31578, -28135, -28666, 
    -23969, -19986, -18817, -14670, -11482, -4847, -2159, 3333, 6955, 11939, 
    13924, 19092, 23056, 24858, 26333, 29719, 31044, 31345, 31525, 31245, 
    28796, 27793, 23197, 20820, 19722, 14019, 11918, 5321, 1567, -1792, 
    -7190, -10936, -15107, -18925, -22002, -26046, -26427, -29791, -30004, 
    -31297, -31911, -29356, -30240, -27409, -25394, -22492, -16987, -15177, 
    -10825, -5638, -2111, 2697, 5729, 11159, 13537, 20155, 22457, 25210, 
    26061, 28221, 30491, 30728, 29582, 30483, 29160, 27018, 24129, 22479, 
    18653, 13717, 10539, 6633, 993, -1798, -6390, -9783, -14572, -17809, 
    -21862, -23737, -26702, -29248, -30009, -30621, -30411, -30815, -28964, 
    -26410, -25016, -23866, -17958, -15330, -10038, -7337, -1725, 2367, 5777, 
    10407, 15247, 17765, 21001, 23294, 26787, 29757, 30708, 29227, 30494, 
    29912, 28616, 27125, 24463, 21251, 19698, 16552, 12409, 6478, 2225, -192, 
    -6268, -9673, -14675, -17364, -20516, -23180, -27598, -27935, -29389, 
    -30273, -30714, -30127, -29147, -27173, -25190, -22153, -19622, -15365, 
    -10743, -6318, -2320, 1385, 5791, 9349, 14133, 16515, 19715, 25214, 
    28090, 27902, 29788, 30838, 31373, 30998, 29205, 27767, 25956, 22562, 
    20661, 16089, 12108, 6896, 2784, -1037, -5501, -9075, -13727, -18111, 
    -20751, -23881, -26094, -28959, -29856, -30839, -30815, -30834, -27718, 
    -27047, -26795, -22606, -19638, -16237, -12265, -8363, -5359, 491, 5171, 
    9158, 12053, 16849, 20198, 23751, 27195, 29077, 29659, 30340, 29020, 
    29569, 29859, 28842, 25802, 22780, 20465, 17056, 12391, 8640, 3130, -412, 
    -3710, -8247, -13550, -16255, -22306, -24240, -25728, -27471, -28527, 
    -29395, -31038, -31219, -29532, -27651, -25408, -22536, -19099, -15896, 
    -11184, -7204, -3979, 499, 4945, 9194, 12973, 17812, 20196, 22724, 26466, 
    28566, 30210, 30388, 31805, 29255, 28790, 26690, 27020, 23143, 20102, 
    16474, 13687, 8083, 4185, -899, -5657, -9894, -13693, -15723, -19748, 
    -23657, -26450, -28067, -28889, -30828, -31168, -31491, -28705, -28234, 
    -25431, -23893, -18955, -15768, -13044, -8261, -4174, 185, 4335, 9013, 
    11990, 15421, 18425, 23961, 26791, 26880, 28750, 30896, 32145, 31119, 
    29273, 27278, 25060, 23767, 21114, 15393, 12846, 9201, 4376, -1313, 
    -4514, -6707, -11963, -17425, -18300, -23194, -24658, -27725, -28952, 
    -30530, -30008, -29837, -29310, -27306, -25568, -22962, -20767, -18021, 
    -13454, -8158, -5661, -477, 2645, 7973, 13033, 16118, 20835, 21525, 
    26331, 28119, 30665, 31530, 31015, 30575, 29411, 27822, 24998, 22985, 
    19726, 18483, 13046, 9811, 3966, 1439, -4500, -8241, -11282, -14793, 
    -21015, -22824, -25404, -26408, -29298, -30590, -31258, -30612, -29636, 
    -28632, -26145, -23915, -20211, -17446, -14643, -9711, -4572, 483, 2618, 
    8207, 11064, 16655, 19191, 22705, 24595, 28161, 30423, 31807, 30843, 
    31304, 28863, 28998, 25213, 23990, 19915, 17587, 13799, 8674, 6941, 284, 
    -3206, -8061, -11458, -15087, -20311, -21107, -25899, -28441, -29982, 
    -29268, -30438, -31609, -30252, -28281, -27230, -23646, -20474, -19142, 
    -13373, -10182, -4460, -408, 3592, 7425, 12699, 16590, 19689, 21838, 
    26043, 27595, 29008, 28720, 31830, 31496, 29313, 29203, 25849, 23487, 
    20728, 19496, 14054, 10208, 6881, 2339, -1589, -7695, -11188, -14538, 
    -19157, -23134, -24815, -26896, -27899, -30406, -29511, -29349, -30884, 
    -27427, -25263, -24360, -22832, -19721, -14573, -11421, -4419, -2531, 
    1939, 6757, 11620, 14693, 18619, 22255, 23771, 28651, 29506, 29457, 
    29711, 30955, 28580, 28020, 27065, 23193, 20618, 18809, 14822, 11179, 
    7322, 2286, -862, -6123, -12465, -14790, -17766, -21748, -24254, -27322, 
    -28245, -29980, -30618, -30651, -29743, -28143, -25741, -25205, -21582, 
    -18159, -16334, -11032, -5217, -1824, 2673, 6459, 12086, 14628, 18357, 
    20813, 25445, 25795, 28323, 28642, 30537, 31920, 29801, 29209, 26806, 
    25290, 21284, 18917, 13552, 12218, 6648, 1869, -3753, -7240, -9939, 
    -14572, -18236, -20054, -24461, -27261, -29263, -28417, -30282, -31678, 
    -31094, -29678, -27229, -24161, -20869, -19382, -16752, -11536, -8119, 
    -3581, 1442, 6953, 11168, 14573, 17594, 23021, 24358, 26950, 27274, 
    29784, 31918, 31595, 28764, 29617, 27803, 25454, 23241, 17478, 15499, 
    11319, 5811, 3657, -709, -6404, -9920, -13496, -18058, -21392, -22891, 
    -27343, -28845, -29789, -29672, -30479, -30002, -29112, -27234, -24281, 
    -22810, -20809, -15434, -10569, -8379, -2692, 989, 7461, 11567, 13856, 
    18584, 20779, 24400, 25619, 27718, 29324, 30989, 31711, 31834, 28962, 
    28534, 24850, 20931, 18667, 15455, 12433, 7816, 2378, -1272, -6644, 
    -9024, -12480, -17671, -21720, -23487, -25388, -27738, -29839, -31712, 
    -30324, -30589, -30268, -26624, -24846, -21964, -20794, -15484, -11025, 
    -6698, -3255, -60, 4121, 10643, 13277, 18355, 22091, 23741, 26969, 28073, 
    29337, 29961, 30093, 30639, 29429, 29255, 24122, 24537, 21566, 15931, 
    12166, 6970, 4908, 118, -4249, -8338, -12696, -16886, -19996, -25071, 
    -26526, -29339, -29743, -30949, -31849, -29817, -27854, -26761, -26667, 
    -23586, -19751, -16265, -12213, -7573, -3675, 521, 5135, 10327, 12998, 
    16916, 20029, 23278, 24825, 28633, 30333, 31458, 29237, 30690, 28942, 
    27822, 24678, 23000, 21718, 17627, 13236, 8768, 5085, -444, -5945, 
    -10517, -13059, -17588, -19305, -23810, -26611, -28331, -28997, -29121, 
    -29580, -30882, -28992, -27116, -26150, -23524, -19848, -18293, -13206, 
    -8404, -3638, 266, 4600, 9059, 11883, 17214, 21501, 24911, 26755, 28125, 
    29367, 31425, 30809, 30942, 29498, 28647, 27569, 22377, 19934, 17208, 
    14082, 10405, 4680, 1343, -3792, -7713, -12103, -15280, -18773, -23953, 
    -27194, -27007, -30441, -29880, -32271, -31848, -30559, -27255, -25444, 
    -23556, -21282, -16984, -12743, -10484, -5729, 714, 4466, 8789, 12200, 
    16840, 19120, 21505, 26232, 27544, 29370, 29036, 29633, 30049, 29471, 
    27811, 26019, 23428, 18981, 16248, 13571, 9970, 4726, 232, -3042, -8809, 
    -12267, -16388, -19564, -21852, -25741, -26802, -30217, -30078, -29291, 
    -30308, -28095, -27372, -25543, -23913, -20985, -18223, -13540, -9070, 
    -5888, 62, 4862, 7882, 12158, 14762, 18996, 21415, 26739, 27685, 30470, 
    30309, 30538, 30209, 29032, 28824, 26642, 24008, 21701, 16073, 13254, 
    9306, 6080, 1998, -3851, -8868, -11095, -15213, -17756, -21540, -25747, 
    -28106, -29602, -30990, -31371, -30470, -29106, -27366, -27691, -24045, 
    -21538, -17544, -13468, -11176, -5714, -1029, 3723, 7151, 11569, 15676, 
    19417, 21927, 26551, 26177, 28605, 29823, 31674, 30816, 29254, 28738, 
    27409, 24856, 20888, 17973, 15262, 10578, 5607, 2774, -2905, -5686, 
    -12306, -14154, -19088, -21672, -24050, -26658, -29838, -28644, -32133, 
    -29362, -29879, -28342, -27455, -23895, -23088, -16676, -14697, -11072, 
    -5847, -1926, 3639, 7626, 11211, 16341, 18232, 23092, 26341, 27643, 
    29206, 30844, 30651, 31305, 30728, 29011, 26236, 25162, 21723, 19010, 
    13863, 10374, 5490, 2828, -1349, -5194, -12135, -15239, -19203, -20421, 
    -25795, -27928, -29365, -29903, -30378, -30723, -29760, -28766, -26809, 
    -23684, -21554, -19219, -15857, -10982, -7572, -3026, 2715, 5886, 11664, 
    14774, 17763, 21584, 24639, 26158, 29305, 29979, 30214, 31617, 29750, 
    28445, 27112, 23513, 22888, 17089, 15719, 10861, 6515, 2406, -1563, 
    -7888, -9452, -14102, -19366, -20870, -22985, -27009, -29346, -30156, 
    -29516, -30224, -30349, -28889, -27248, -24213, -22896, -19038, -14393, 
    -11169, -7172, -3393, 478, 6404, 9764, 15055, 17609, 21594, 24466, 26110, 
    28288, 30480, 29809, 30192, 29583, 29180, 26353, 24146, 20536, 19404, 
    16876, 10973, 6669, 2896, -2469, -5485, -10550, -15825, -17395, -21339, 
    -24056, -25886, -28008, -30366, -31661, -30340, -29342, -27877, -27286, 
    -23748, -22879, -20216, -15224, -10228, -6291, -2726, -603, 6205, 10083, 
    14168, 16661, 21907, 23934, 27559, 28460, 29821, 30276, 31220, 29831, 
    30613, 27475, 25247, 23430, 19322, 16201, 10749, 9006, 1675, -1152, 
    -7194, -9139, -12379, -18521, -21752, -23659, -25978, -29051, -29355, 
    -32208, -30429, -30419, -29191, -28210, -25105, -24232, -20593, -14644, 
    -11688, -7244, -1899, 2055, 4290, 8738, 13620, 18522, 20000, 23861, 
    24747, 27352, 30090, 32222, 31963, 30893, 30536, 26469, 26206, 22889, 
    19410, 16676, 13227, 7623, 3973, 1137, -4300, -9603, -14992, -17580, 
    -20762, -23489, -26944, -27257, -28207, -30455, -30913, -30297, -28991, 
    -26717, -25741, -23223, -19089, -15787, -11661, -8811, -3986, 53, 4740, 
    9738, 15016, 17006, 21444, 23219, 25491, 28967, 28473, 30030, 30965, 
    32094, 29728, 27650, 24630, 22505, 19004, 16476, 12259, 8153, 3146, 279, 
    -5193, -9910, -13129, -16662, -21142, -22486, -26027, -27594, -29347, 
    -30973, -30160, -31523, -28310, -27477, -25810, -23908, -19639, -17378, 
    -14203, -8342, -4086, -658, 5755, 7808, 13206, 16134, 19722, 23838, 
    27308, 27337, 28625, 30643, 31900, 31281, 28244, 27963, 24589, 24620, 
    20721, 17075, 12853, 8874, 5168, -198, -4803, -8345, -11710, -16058, 
    -20117, -23076, -25605, -27899, -30281, -29933, -31583, -30497, -30190, 
    -27003, -27007, -23730, -20072, -16579, -12165, -8252, -4938, 379, 3726, 
    7667, 14236, 14670, 20216, 22940, 26143, 28464, 30178, 31028, 31371, 
    31692, 29038, 27971, 24883, 22132, 20937, 17239, 12202, 10529, 4055, 
    1491, -3098, -8769, -12450, -15388, -19605, -24298, -25720, -29248, 
    -29452, -31065, -31771, -29301, -29529, -27202, -26032, -24851, -20890, 
    -18129, -13224, -9375, -5770, -818, 2664, 7818, 11958, 15411, 19033, 
    22697, 24564, 27076, 29429, 30179, 31500, 30862, 29389, 28781, 26298, 
    22870, 21164, 18208, 13231, 8114, 5378, -620, -4661, -6952, -11241, 
    -15238, -17526, -21231, -24847, -27364, -28728, -29054, -30503, -30521, 
    -30619, -28000, -28027, -22667, -20946, -18733, -13948, -10652, -5271, 
    -458, 1776, 7189, 10840, 16541, 18267, 23743, 25888, 27590, 29250, 28937, 
    30660, 30419, 31326, 28484, 26697, 24895, 19496, 16724, 14347, 9436, 
    6536, 480, -3179, -6522, -9587, -15370, -19017, -22428, -25047, -27870, 
    -30536, -30366, -29573, -30609, -30169, -28240, -25454, -23952, -21382, 
    -17194, -15137, -9296, -6983, -492, 1963, 7394, 11331, 14113, 19387, 
    22098, 25891, 27672, 29077, 29339, 31188, 31776, 30148, 27801, 27297, 
    24338, 21018, 18954, 14255, 10402, 5705, 2271, -3350, -8198, -11046, 
    -15383, -18988, -21150, -23986, -26999, -29633, -29847, -32111, -29287, 
    -30009, -29008, -26105, -24663, -22261, -19176, -14339, -11159, -5740, 
    -1258, 2142, 6729, 10304, 15744, 18095, 21144, 25376, 26574, 28036, 
    29596, 31094, 31367, 31629, 27503, 26779, 24721, 22446, 18951, 14338, 
    10646, 6414, 2727, -2470, -5348, -12254, -13911, -18196, -21545, -24951, 
    -27810, -28710, -30566, -30724, -31651, -30798, -27721, -27135, -25181, 
    -21649, -19171, -16347, -10496, -7625, -2383, 903, 5362, 10732, 14939, 
    18130, 21731, 24790, 25209, 29501, 30239, 30808, 30901, 29875, 29205, 
    26610, 24388, 21558, 19371, 14735, 11170, 6064, 4042, -1654, -5292, 
    -10030, -14125, -18448, -20589, -24012, -27710, -29211, -29161, -31110, 
    -31340, -32085, -30209, -26536, -24651, -22955, -17902, -15015, -11023, 
    -7683, -4144, 1547, 4181, 9494, 13507, 17364, 21542, 24180, 27683, 29637, 
    30063, 31680, 29694, 31319, 29860, 28055, 26793, 22264, 20621, 15742, 
    11509, 9262, 2260, -45, -6376, -8953, -14186, -16304, -19673, -24893, 
    -25920, -28449, -30834, -31437, -31099, -28932, -30217, -27306, -25508, 
    -21359, -20795, -16394, -12487, -6961, -3525, 1131, 5128, 8018, 14356, 
    16761, 19775, 24608, 26791, 26829, 31311, 30102, 30057, 31601, 29362, 
    28752, 25026, 21656, 19234, 14854, 12240, 7600, 3626, -1181, -4721, 
    -8043, -13736, -16757, -21118, -23223, -25577, -28891, -29833, -29463, 
    -30812, -30452, -30242, -28514, -26850, -21839, -19439, -17632, -11300, 
    -8662, -4343, 369, 5184, 8829, 13807, 17161, 21347, 23238, 25972, 28677, 
    28811, 30590, 32545, 30822, 29902, 28486, 24717, 23841, 21307, 14979, 
    11164, 7556, 5463, -418, -5302, -7361, -11144, -16246, -19367, -22371, 
    -24678, -28487, -29291, -30083, -31544, -30194, -29777, -28498, -26063, 
    -22701, -20177, -15526, -11415, -8968, -4520, -538, 3503, 7745, 12812, 
    17533, 21185, 23503, 25756, 29363, 29736, 29204, 30662, 30838, 30925, 
    26720, 27608, 24086, 18523, 16626, 12614, 9299, 5739, -12, -4392, -7337, 
    -12900, -17293, -19843, -22561, -24982, -28975, -28540, -32033, -32320, 
    -31461, -29615, -28553, -24818, -22912, -20704, -17503, -14287, -9720, 
    -3323, -736, 4156, 8871, 12208, 16648, 19114, 23388, 25325, 29272, 28162, 
    29546, 30391, 30100, 29470, 27403, 26271, 23593, 20061, 17361, 12959, 
    10312, 4341, 537, -3571, -8564, -10464, -16403, -19456, -22142, -25875, 
    -27179, -30291, -30598, -31251, -30350, -28861, -29330, -25834, -24082, 
    -22147, -18098, -13191, -10196, -5151, -1924, 2845, 8054, 11311, 16162, 
    20670, 22685, 25483, 26952, 29699, 31055, 30332, 29687, 29703, 27748, 
    27513, 24359, 19858, 16630, 14767, 8473, 5839, 60, -2849, -8204, -12025, 
    -15759, -18653, -23197, -24514, -26228, -28928, -30536, -31053, -30381, 
    -30201, -27739, -26246, -23229, -22171, -16725, -13338, -11045, -4409, 
    -2318, 4228, 8861, 11886, 15498, 19917, 21965, 23398, 28033, 30894, 
    30413, 32487, 31080, 30613, 27917, 26690, 23539, 21725, 16196, 13282, 
    10540, 6177, 544, -3999, -8532, -10579, -15990, -18443, -22143, -26229, 
    -27831, -28384, -30336, -31433, -30370, -30097, -29853, -27003, -23517, 
    -22216, -18475, -13554, -10934, -5842, -2776, 3774, 6990, 11916, 15914, 
    18730, 21083, 24335, 28433, 29280, 30248, 31138, 31483, 30699, 28525, 
    28208, 24815, 23140, 18146, 15436, 10950, 6137, 1736, -2692, -6538, 
    -10836, -15241, -19830, -22144, -24254, -28922, -29453, -30274, -29757, 
    -32290, -30876, -29341, -27200, -26024, -21563, -17856, -15691, -11455, 
    -6472, -1736, 2173, 7224, 10517, 14383, 18351, 21070, 25700, 28152, 
    29043, 31801, 30436, 30366, 30235, 27699, 28573, 24026, 21876, 18542, 
    13705, 10985, 6786, 3044, -2523, -7333, -9948, -14565, -17905, -20774, 
    -24691, -26564, -29208, -29304, -29940, -30104, -29951, -29129, -26686, 
    -23977, -21646, -18054, -15080, -10844, -7187, -2321, 1770, 4928, 10460, 
    14491, 18263, 21657, 23916, 27105, 28702, 29047, 32319, 31572, 31102, 
    29281, 26203, 25387, 22162, 19986, 15811, 12144, 8331, 3006, -2298, 
    -6953, -9824, -14073, -17807, -21489, -25294, -27219, -28728, -30205, 
    -30493, -32178, -28980, -28576, -27188, -24657, -23069, -19545, -16719, 
    -9867, -7323, -2404, 2503, 5921, 10469, 13505, 18442, 20266, 24707, 
    26285, 27741, 29548, 29781, 29449, 30308, 31124, 28778, 26148, 22850, 
    18482, 15645, 11016, 8511, 4101, -1305, -4780, -10483, -13479, -16177, 
    -22244, -23892, -25426, -27638, -29667, -30492, -31685, -29907, -30562, 
    -28113, -25139, -23076, -18935, -15044, -12354, -7503, -2684, 1261, 5057, 
    10633, 14238, 17262, 22162, 23733, 26503, 28881, 30103, 30769, 31385, 
    30502, 30394, 27083, 26025, 22589, 18914, 16192, 11128, 6300, 5414, 
    -1179, -4814, -7814, -13106, -16159, -20152, -23425, -25702, -26988, 
    -30239, -30260, -31918, -31480, -29631, -26720, -25472, -23274, -19932, 
    -14988, -12595, -7127, -3577, 459, 5120, 9581, 13095, 16654, 19028, 
    23668, 24701, 28186, 30809, 29094, 31294, 30579, 30322, 28612, 26410, 
    22576, 18987, 16956, 12943, 9042, 4535, -485, -5755, -9266, -13456, 
    -17586, -20530, -23831, -26078, -26718, -31385, -30532, -31272, -30154, 
    -29769, -28481, -24826, -24194, -19547, -16589, -12406, -8185, -4513, 
    575, 6095, 8920, 12903, 17086, 19532, 23605, 25318, 28023, 29168, 29297, 
    31175, 31351, 28983, 26548, 27189, 22995, 19859, 16479, 13078, 7978, 
    4805, 498, -5179, -9261, -11356, -17410, -21144, -24181, -27361, -27542, 
    -28805, -30221, -32035, -31175, -29628, -28784, -25919, -22316, -21990, 
    -17606, -13404, -7898, -5708, -1948, 5614, 7481, 11943, 17904, 19157, 
    23486, 23982, 28140, 29280, 30192, 31121, 30997, 28980, 28502, 26924, 
    24774, 20749, 16300, 12773, 9673, 4580, 363, -4193, -7795, -12160, 
    -16411, -18336, -21377, -25424, -27466, -29779, -30452, -30232, -29091, 
    -29622, -28175, -26309, -25043, -21945, -18523, -13630, -9328, -6486, 
    -1766, 4723, 8687, 11906, 15177, 20075, 24182, 25670, 27939, 29175, 
    31277, 30478, 31703, 29118, 28409, 26456, 23127, 20848, 16654, 14197, 
    8627, 5441, 489, -4819, -8207, -11333, -14766, -19447, -22946, -25320, 
    -26568, -28196, -29393, -31211, -31466, -29789, -28625, -25733, -25359, 
    -21385, -18359, -14427, -11093, -6069, -1302, 1542, 8000, 11782, 16637, 
    19441, 21258, 25474, 28242, 29010, 30847, 30482, 30264, 31178, 28469, 
    26183, 23892, 22656, 17529, 14322, 9956, 6320, 790, -3960, -5658, -11489, 
    -15841, -18828, -21465, -24832, -28386, -28647, -31169, -30749, -30631, 
    -30066, -28357, -26154, -23630, -19657, -18716, -14139, -11186, -6770, 
    -2666, 1890, 7076, 10980, 15244, 18579, 21567, 23865, 28701, 27142, 
    29481, 30558, 31512, 30635, 27563, 26757, 24410, 21265, 17272, 13875, 
    8814, 4916, 2682, -1460, -7239, -10790, -14956, -19009, -21934, -25675, 
    -28176, -28255, -29992, -31616, -32272, -29134, -28813, -28397, -24602, 
    -21536, -18601, -14008, -9329, -6034, -1987, 2247, 8019, 9994, 14786, 
    18079, 22430, 25918, 26659, 29323, 29152, 29986, 30193, 30207, 28617, 
    27319, 25035, 22282, 18506, 14132, 10144, 6390, 3820, -887, -5884, 
    -11242, -15821, -19323, -22990, -23832, -26932, -28127, -29757, -29524, 
    -30092, -29558, -28515, -27346, -25175, -22462, -17510, -14812, -9804, 
    -8374, -1731, 3307, 7136, 10616, 14159, 18240, 21429, 24500, 27185, 
    28237, 29885, 31005, 31182, 31571, 29929, 27169, 24576, 22345, 17995, 
    15167, 12963, 6318, 4007, -3007, -5334, -10005, -14425, -16700, -19998, 
    -23694, -26440, -27826, -29161, -30671, -31484, -29816, -29049, -27041, 
    -24063, -23403, -18994, -15932, -11179, -8661, -4055, 1671, 5707, 9812, 
    12545, 19011, 21832, 23791, 27359, 29212, 29851, 29780, 30383, 30434, 
    29620, 28869, 25004, 22206, 19361, 15572, 13602, 8134, 4788, -1712, 
    -4738, -10600, -12566, -16623, -20271, -23513, -26787, -28081, -30605, 
    -30886, -31215, -30420, -29888, -27129, -26066, -22875, -19170, -14928, 
    -12068, -8934, -4673, 495, 6657, 10602, 14102, 17537, 20041, 23444, 
    25336, 28790, 28828, 30209, 32047, 30598, 29601, 27271, 25935, 23761, 
    18086, 15563, 12330, 8992, 2707, -1791, -5151, -9362, -14382, -17396, 
    -19917, -22757, -24329, -28163, -30163, -30265, -30307, -30804, -29545, 
    -27281, -25494, -23071, -20970, -17284, -11529, -8481, -4678, 214, 4911, 
    9149, 12744, 16841, 19738, 23653, 25038, 27807, 29264, 31970, 30631, 
    30295, 29322, 27206, 26399, 22722, 21034, 17666, 13694, 8475, 3488, -276, 
    -4841, -9564, -13631, -16257, -20049, -24082, -25720, -27628, -29405, 
    -30766, -30124, -30583, -29127, -28202, -25033, -22856, -19741, -17513, 
    -13853, -9958, -5352, 433, 4482, 8555, 11390, 16550, 20323, 23880, 26754, 
    26485, 29050, 29747, 31036, 29443, 28775, 27642, 26145, 24116, 20774, 
    17192, 14663, 9025, 4619, 639, -2839, -6902, -12566, -17928, -20135, 
    -22213, -25466, -28553, -30224, -30442, -30841, -31291, -28622, -27310, 
    -25949, -22915, -20408, -17673, -12464, -10446, -5443, -603, 2028, 8856, 
    11615, 16758, 20378, 23054, 26981, 28758, 29380, 29459, 29487, 30560, 
    30992, 28690, 26432, 24268, 19943, 15564, 13714, 10076, 4653, -361, 
    -4962, -6533, -12147, -16439, -19637, -22448, -24820, -28537, -28197, 
    -29796, -32338, -30861, -29485, -28495, -26555, -25560, -20161, -17189, 
    -15083, -8548, -4703, -1190, 2947, 6249, 12495, 17455, 18718, 21235, 
    25531, 28627, 28512, 30971, 30865, 31437, 28518, 28392, 26472, 23373, 
    20148, 17587, 13572, 9451, 4263, -140, -3069, -7579, -12451, -16316, 
    -18164, -22726, -25853, -27778, -27819, -30857, -31697, -30203, -29971, 
    -29054, -27006, -25290, -20756, -18749, -15016, -10011, -4083, -1557, 
    3984, 7376, 10937, 15602, 18838, 22717, 26349, 27114, 28636, 29747, 
    30558, 30926, 30211, 28765, 27138, 24021, 22051, 18539, 13758, 10144, 
    6791, 2302, -3422, -7541, -11617, -15366, -18078, -21451, -24115, -26955, 
    -29061, -30904, -30899, -32542, -28668, -28469, -26774, -23186, -21894, 
    -17171, -13407, -10535, -6372, -1972, 2520, 8152, 11224, 15272, 19282, 
    21167, 24220, 27363, 30611, 29674, 30813, 30337, 29250, 29661, 26439, 
    23342, 21061, 17953, 14303, 11018, 6677, 2628, -3032, -7208, -11120, 
    -15180, -17863, -21902, -25056, -27502, -29968, -30296, -31405, -31545, 
    -30527, -27983, -26527, -24265, -22833, -17896, -14795, -12085, -7612, 
    -1325, 3456, 5122, 10756, 15942, 17095, 23147, 24041, 27298, 28212, 
    30153, 29400, 30505, 30900, 28008, 28083, 24167, 21995, 17414, 15096, 
    10661, 6539, 1063, -3443, -6324, -9863, -14611, -17619, -21596, -25987, 
    -26554, -29741, -31045, -31157, -31056, -30001, -28687, -28543, -23700, 
    -22558, -19080, -15381, -12497, -6510, -2037, 2295, 6364, 8633, 13917, 
    18624, 22552, 22671, 27367, 29101, 30171, 31097, 30251, 29283, 30148, 
    28208, 24274, 22140, 19758, 16703, 12676, 6547, 2125, -1655, -5589, 
    -10424, -15414, -17307, -19626, -25715, -25977, -28421, -30071, -29865, 
    -30312, -29688, -28172, -27873, -26522, -22386, -19391, -15094, -13050, 
    -6544, -3786, 739, 4952, 9861, 12960, 18663, 21224, 23344, 26106, 28656, 
    29966, 31494, 30254, 30267, 28713, 28802, 26551, 21052, 20051, 14834, 
    11070, 6942, 4116, -991, -5227, -10220, -12807, -17382, -20579, -23013, 
    -26354, -28993, -28476, -30846, -31041, -30291, -29318, -27343, -25090, 
    -23206, -20503, -14601, -12929, -8842, -3552, 477, 4428, 9631, 15022, 
    18054, 19915, 24332, 24962, 28032, 28298, 31402, 32506, 29209, 29547, 
    27343, 25349, 22090, 19389, 15736, 12059, 8105, 3704, -1056, -6024, 
    -8735, -11809, -16062, -19533, -23342, -27256, -28329, -29648, -29810, 
    -31433, -30782, -28198, -27755, -25600, -23222, -20326, -16693, -11939, 
    -7482, -3932, 334, 4897, 8220, 12426, 17421, 20419, 22650, 24849, 28403, 
    28977, 31345, 31522, 30944, 27611, 27321, 25380, 23744, 20722, 16109, 
    12663, 8209, 3886, 151, -4987, -9376, -12939, -16770, -20558, -22746, 
    -26087, -28038, -30066, -31266, -30311, -31000, -29665, -28296, -26526, 
    -23956, -20343, -16485, -11761, -8625, -4418, 712, 4206, 9852, 12588, 
    16290, 19467, 23142, 26088, 28612, 29389, 31383, 32270, 32369, 30980, 
    28840, 27106, 22135, 20304, 17499, 13754, 8144, 3991, 1697, -5115, -8227, 
    -13964, -16650, -20734, -23322, -25169, -28321, -30051, -30494, -29854, 
    -30849, -30391, -29373, -26675, -23113, -19829, -17382, -13831, -9285, 
    -4870, -209, 2517, 7463, 11754, 17535, 19604, 21772, 25952, 28162, 29921, 
    30469, 30695, 29816, 29959, 26501, 27162, 22765, 21986, 16919, 13230, 
    8206, 4726, 535, -2315, -6604, -12136, -14982, -19910, -21970, -25709, 
    -26195, -29418, -29009, -31028, -29979, -29608, -28172, -25954, -23512, 
    -20267, -18353, -13764, -9657, -5540, -1062, 2487, 7807, 12908, 15783, 
    20155, 23450, 25408, 27771, 29322, 31135, 30676, 29801, 29817, 28189, 
    28048, 24546, 21856, 16387, 14223, 10098, 4983, 1506, -3925, -6615, 
    -10797, -16280, -19289, -22945, -24210, -27797, -29486, -29138, -29495, 
    -29894, -30612, -28300, -26642, -24972, -20536, -19227, -13826, -10364, 
    -5674, -116, 3172, 7479, 12142, 16453, 19373, 22423, 25674, 27512, 29242, 
    30101, 31350, 30169, 30590, 28671, 27855, 24745, 21563, 18388, 13385, 
    10711, 5912, -288, -3003, -7176, -12854, -14415, -18563, -23701, -24901, 
    -26215, -29707, -29090, -31451, -30713, -31080, -28526, -27358, -22554, 
    -20353, -16707, -14449, -10188, -4524, -2502, 3123, 7320, 11726, 15420, 
    18030, 23005, 24288, 28344, 30563, 29753, 31436, 31815, 29706, 27397, 
    27055, 25368, 21712, 18907, 13968, 10923, 4810, 3169, -1684, -6390, 
    -10884, -14154, -17421, -20631, -23505, -26427, -28692, -30170, -31085, 
    -30379, -29442, -29511, -27235, -24697, -22264, -18392, -14046, -12083, 
    -4791, -697, 1072, 6910, 11301, 15111, 18645, 20942, 24298, 25383, 29222, 
    29736, 29191, 32457, 29949, 28351, 26963, 25469, 20599, 17465, 15088, 
    10353, 7953, 2527, -2015, -6310, -10721, -14343, -17521, -21153, -24539, 
    -26036, -29591, -28916, -31263, -32103, -29785, -29363, -26692, -25204, 
    -22462, -18413, -15136, -10207, -6848, -4091, 1970, 6342, 10280, 12952, 
    18397, 21222, 23515, 25965, 27093, 31630, 29657, 29616, 29461, 27708, 
    25829, 24617, 22186, 18894, 14113, 11307, 6003, 2472, -1117, -6562, 
    -10873, -14849, -19156, -21273, -24106, -27576, -28497, -29188, -29745, 
    -30927, -29746, -29388, -26758, -26248, -23464, -20184, -15379, -10503, 
    -7322, -2945, 1137, 5567, 9742, 14526, 17090, 20421, 24688, 26382, 28784, 
    29561, 31973, 30903, 30686, 28277, 28018, 25900, 22207, 19082, 14381, 
    10597, 7253, 2136, -2426, -4252, -9601, -14321, -16425, -20577, -24269, 
    -26058, -28557, -31389, -31108, -29929, -30279, -28666, -26925, -24933, 
    -23952, -18840, -16636, -10950, -7890, -2829, -956, 5211, 9951, 15210, 
    18816, 21602, 23776, 25097, 28228, 29464, 29825, 30766, 29382, 28136, 
    27436, 24815, 22940, 19377, 14963, 12255, 8188, 2208, -184, -4110, -8610, 
    -14230, -18176, -20208, -24607, -26135, -29352, -29966, -30052, -31647, 
    -30354, -30786, -27383, -25606, -24642, -19137, -16983, -13381, -7055, 
    -3153, 48, 4930, 9345, 14337, 17563, 21498, 23043, 25722, 27833, 28997, 
    30828, 31469, 30377, 28245, 27411, 26843, 24175, 19139, 17408, 12552, 
    8258, 3799, 600, -5771, -9451, -13703, -16959, -19393, -23948, -24780, 
    -26435, -28880, -30140, -29974, -29923, -29678, -27851, -25451, -22999, 
    -18858, -16825, -12482, -7978, -3411, 936, 3264, 8861, 13316, 17345, 
    20568, 22253, 25915, 27993, 30006, 30738, 32468, 29784, 29847, 27057, 
    25658, 23413, 21404, 18420, 13657, 8603, 4878, 614, -3221, -8469, -12584, 
    -16761, -20221, -22610, -25542, -28885, -28421, -30000, -29775, -29471, 
    -30901, -28830, -25831, -23963, -19905, -15807, -12477, -9287, -6030, 
    346, 4740, 8000, 11357, 16856, 18932, 22999, 27196, 27759, 29124, 29912, 
    30979, 29777, 29456, 28487, 25551, 23347, 20557, 15633, 11587, 8388, 
    5934, 873, -4144, -7773, -11144, -14590, -19311, -23171, -26081, -26792, 
    -29966, -31383, -30039, -32012, -30697, -29477, -26619, -23958, -20466, 
    -17930, -13203, -9976, -6073, -67, 3197, 8191, 12322, 14993, 19608, 
    22836, 24789, 28942, 29275, 29879, 29821, 31496, 30813, 28045, 26442, 
    23314, 20643, 18753, 14738, 10324, 5430, 698, -3134, -7272, -10226, 
    -15585, -19396, -22010, -25622, -27256, -29619, -30227, -30848, -30013, 
    -30477, -29822, -26864, -22607, -21229, -17770, -14168, -8972, -4787, 
    -764, 3483, 5930, 11710, 15928, 19594, 22507, 24245, 26088, 29291, 29395, 
    31187, 29420, 29194, 28403, 25908, 23869, 22072, 19377, 15298, 10189, 
    4499, 1098, -2027, -6907, -11906, -15571, -18070, -22723, -25130, -28683, 
    -27824, -31517, -29177, -29735, -30428, -29609, -27855, -23260, -22424, 
    -18259, -15198, -11009, -6110, -2191, 3784, 6841, 12261, 16183, 17979, 
    21056, 24489, 27097, 28606, 29741, 31850, 30507, 30179, 28791, 26539, 
    25041, 21461, 18644, 14581, 9166, 7264, 1802, -1554, -7414, -10915, 
    -13244, -18407, -22795, -24060, -26662, -29795, -29653, -30718, -31353, 
    -29451, -27606, -26987, -26234, -21284, -17837, -15636, -11607, -5913, 
    -3122, 2762, 8121, 11891, 14540, 17689, 22087, 25691, 26682, 27583, 
    29828, 29564, 30105, 29078, 30305, 25326, 24092, 20690, 17479, 14849, 
    10158, 7068, 3630, -3221, -5766, -11806, -15084, -18672, -22155, -23453, 
    -28102, -28909, -30122, -31097, -30955, -31379, -29184, -27641, -26428, 
    -21708, -17566, -15971, -11705, -6986, -3385, 353, 5796, 10575, 13704, 
    17092, 20118, 24952, 27967, 29286, 28577, 28965, 30122, 30694, 29048, 
    27835, 26410, 23824, 19940, 16472, 11661, 7191, 2646, -1929, -4697, 
    -9699, -15473, -18086, -22495, -23674, -26976, -29475, -28878, -30622, 
    -30778, -30349, -29119, -26219, -25042, -21064, -18964, -16045, -11373, 
    -7305, -3159, 1966, 5362, 8960, 15632, 18550, 21430, 23193, 26627, 27161, 
    28758, 31444, 29501, 31659, 28245, 26895, 24809, 21881, 18604, 16545, 
    12828, 8060, 3199, -499, -5193, -8408, -14235, -17230, -21238, -22618, 
    -25272, -27211, -29175, -30068, -32460, -31598, -29846, -28859, -26206, 
    -20797, -20434, -15733, -13764, -6263, -2795, 832, 4727, 10383, 12509, 
    17103, 21670, 23771, 25679, 29169, 30624, 30362, 31717, 31435, 30410, 
    27453, 25003, 23769, 20264, 16739, 12208, 7563, 3322, -1308, -3404, 
    -9931, -13283, -16999, -21539, -24161, -27194, -27159, -29686, -30862, 
    -30768, -30025, -29129, -27771, -26343, -23925, -19954, -16056, -12021, 
    -9459, -3100, 676, 3896, 8806, 12210, 17767, 21838, 22832, 26434, 27009, 
    30914, 29114, 30393, 31190, 29053, 28191, 25867, 22579, 20625, 17059, 
    11826, 8661, 4879, -407, -3563, -8296, -13743, -16094, -19471, -23736, 
    -26101, -27076, -28693, -31823, -31133, -30025, -29572, -28619, -27337, 
    -23303, -20250, -16927, -13635, -8700, -6104, -974, 4422, 9297, 12727, 
    17402, 20465, 22511, 24819, 28987, 29089, 29530, 29415, 30215, 29026, 
    27923, 26451, 23611, 21264, 16895, 13012, 9004, 3811, 424, -4164, -9162, 
    -11635, -16782, -18871, -21619, -24953, -26602, -28743, -30323, -30749, 
    -30837, -29189, -27854, -26855, -23412, -18860, -17334, -12785, -9135, 
    -4671, -820, 4523, 7202, 11146, 17192, 18917, 24204, 24687, 28264, 29266, 
    29530, 31470, 29659, 29496, 29551, 24708, 23314, 20836, 17521, 11731, 
    7587, 3199, 554, -4102, -9101, -11512, -15582, -19497, -21160, -26155, 
    -29125, -30129, -31678, -31250, -29883, -29956, -27453, -26654, -23765, 
    -22042, -15961, -13704, -10227, -5610, -1595, 3386, 9624, 12071, 15160, 
    20380, 21357, 25383, 26997, 28003, 31944, 29983, 31862, 29703, 27989, 
    27418, 22713, 21340, 18290, 12890, 8934, 4486, 1051, -1492, -8389, 
    -11458, -13885, -19248, -21653, -25765, -26628, -30705, -29871, -30491, 
    -30447, -31306, -28781, -25825, -24167, -20270, -18187, -13727, -8600, 
    -4712, -1077, 3086, 7775, 12294, 15740, 18627, 22866, 26315, 26923, 
    28839, 31467, 29729, 29507, 28440, 28722, 26569, 22883, 22255, 18171, 
    14965, 9346, 5958, 876, -2715, -6802, -11864, -15447, -18828, -21426, 
    -25703, -27818, -30050, -31546, -32321, -30434, -29908, -28854, -26184, 
    -24653, -22552, -16316, -14021, -9124, -6949, -2935, 2211, 7203, 12163, 
    15515, 19370, 23502, 25203, 27258, 29120, 28343, 30013, 31200, 30819, 
    28904, 25803, 23799, 21946, 18722, 13608, 9839, 4650, 2311, -2770, -7672, 
    -11109, -16587, -17190, -21407, -25033, -26450, -30250, -29922, -31559, 
    -31043, -29698, -30725, -26485, -23942, -21224, -16957, -15252, -11253, 
    -6359, -2805, 2615, 6951, 10915, 15680, 18326, 20526, 25577, 25987, 
    29689, 29898, 30705, 30216, 29257, 29125, 27478, 26607, 22467, 18848, 
    14485, 11126, 7483, 2279, -1125, -6881, -11438, -14386, -19088, -21394, 
    -23422, -26527, -27433, -29744, -30557, -30365, -29033, -29064, -26843, 
    -26169, -21413, -20306, -15706, -11357, -7229, -4017, 2109, 5483, 9309, 
    14587, 19661, 20067, 24325, 26497, 28506, 30204, 30005, 31038, 28714, 
    29087, 27059, 23729, 22248, 20681, 14515, 11983, 6912, 2630, -2476, 
    -5655, -9770, -15342, -17897, -20727, -25066, -25208, -27129, -29959, 
    -31001, -31091, -29734, -29280, -27794, -24777, -22370, -19319, -15678, 
    -11415, -8837, -2680, 214, 6093, 9820, 13412, 18912, 21651, 24047, 26236, 
    29355, 30085, 29504, 30746, 30608, 28671, 28350, 25430, 21863, 19475, 
    15675, 11039, 6631, 4385, -533, -6359, -10378, -13438, -17745, -19413, 
    -25619, -25377, -29004, -30203, -30041, -29253, -31049, -30190, -27936, 
    -25761, -22613, -20803, -16575, -12608, -8159, -4391, 1537, 4353, 10521, 
    13555, 18519, 21693, 25481, 26264, 28687, 29407, 30970, 30981, 29843, 
    30437, 29134, 25637, 23508, 20182, 16936, 13886, 7940, 3436, -1135, 
    -4897, -8910, -13392, -17304, -19751, -22926, -25354, -27637, -29991, 
    -30579, -30670, -29953, -28574, -27835, -26694, -21676, -18344, -16574, 
    -13297, -6977, -4464, 1144, 4222, 10144, 13566, 17550, 20350, 23319, 
    24770, 29160, 30567, 30729, 31961, 30812, 29976, 27681, 25568, 24145, 
    20541, 17375, 12512, 9197, 5200, -1157, -4965, -7960, -11623, -15403, 
    -20677, -22416, -26600, -27378, -28395, -30584, -30959, -29689, -30011, 
    -28633, -27349, -22342, -20191, -16494, -11387, -7777, -5591, -1393, 
    4513, 8752, 13326, 16520, 20161, 22931, 25643, 27472, 29817, 31025, 
    29875, 31802, 29114, 28779, 25816, 23725, 20856, 16864, 12822, 8689, 
    3805, 983, -3638, -7906, -12694, -17161, -20349, -23543, -26345, -28560, 
    -30059, -30458, -30994, -31306, -31083, -29166, -25248, -23638, -19292, 
    -16458, -12994, -8216, -2962, -2054, 4328, 7944, 11977, 15908, 20282, 
    21607, 27147, 28868, 29482, 31477, 31295, 30280, 31123, 29834, 25667, 
    23192, 19707, 16262, 13098, 8973, 5485, 208, -2715, -7917, -11267, 
    -15317, -19242, -22259, -24326, -27777, -28334, -31119, -31495, -31536, 
    -29251, -29416, -27240, -24051, -22118, -16881, -14386, -9678, -6760, 
    -662, 2137, 8628, 13060, 14135, 19964, 22370, 25622, 28163, 30280, 29764, 
    32113, 29667, 29621, 27872, 25873, 23957, 20831, 17125, 13065, 9037, 
    6789, 2434, -3055, -7456, -11464, -16762, -17872, -21747, -26094, -26432, 
    -27819, -30654, -30035, -30835, -29349, -28612, -26604, -23258, -21630, 
    -16123, -13575, -10741, -4932, -1901, 2198, 8290, 9796, 16782, 19602, 
    22010, 24559, 27178, 28945, 31538, 30989, 31992, 30032, 29954, 27005, 
    24935, 20065, 18996, 14689, 9618, 7298, 977, -3294, -6324, -9767, -17073, 
    -18916, -22272, -25472, -28113, -30424, -31165, -30186, -32225, -31108, 
    -29647, -27249, -24370, -21263, -18279, -14604, -10887, -6103, -3219, 
    2949, 7517, 10664, 14169, 19362, 21990, 23745, 26435, 29004, 30698, 
    32572, 30075, 29736, 30020, 27367, 22981, 20989, 18136, 14730, 10224, 
    6289, 2993, -2917, -7138, -11485, -14407, -18150, -21215, -26319, -28684, 
    -27766, -30554, -29805, -28952, -30783, -28439, -27618, -24986, -22439, 
    -20116, -14857, -10772, -7198, -706, 500, 6310, 10078, 12905, 17288, 
    21335, 25407, 26084, 29684, 29997, 30825, 30326, 30781, 28073, 26206, 
    24516, 20895, 19387, 16224, 9589, 6710, 999, -1940, -6629, -10741, 
    -14165, -17237, -21383, -24003, -26280, -29035, -30346, -31133, -31493, 
    -31039, -29034, -28375, -26222, -22317, -19871, -14193, -11073, -6237, 
    -3231, 3286, 5726, 11058, 14466, 18641, 22675, 24331, 26355, 27917, 
    30066, 30712, 30334, 30726, 29370, 28426, 23605, 21567, 18391, 16183, 
    11445, 6980, 4169, -1083, -6866, -11786, -14693, -19530, -20370, -24279, 
    -25972, -27144, -28433, -30055, -30917, -29950, -30045, -26996, -24752, 
    -23685, -18742, -14882, -11790, -7843, -4296, -432, 5172, 10490, 12703, 
    17490, 22232, 24695, 27490, 27663, 29607, 30548, 29039, 30490, 27641, 
    27394, 24268, 22053, 18310, 16110, 12341, 7889, 3065, -474, -5583, -9959, 
    -12932, -16630, -21771, -23761, -25487, -29507, -29831, -29121, -30757, 
    -29889, -29078, -26429, -24737, -23933, -20945, -16186, -12068, -7873, 
    -2984, 295, 5034, 9159, 12285, 16718, 22659, 23392, 25345, 29281, 28994, 
    31056, 30564, 30055, 28595, 28110, 25376, 22643, 20783, 16491, 12281, 
    9247, 3845, -793, -4477, -8150, -12469, -18199, -19684, -23956, -24714, 
    -29063, -28730, -29719, -30783, -29468, -29575, -26764, -25014, -22036, 
    -18685, -17191, -12404, -7663, -2065, -197, 4915, 9638, 13572, 16433, 
    20100, 23945, 25909, 28158, 29500, 30347, 30086, 31459, 30197, 27112, 
    26424, 22504, 18362, 14674, 13220, 9988, 5620, 938, -4407, -8445, -12655, 
    -16164, -20614, -22427, -26008, -28233, -29925, -30515, -30681, -31451, 
    -30659, -27105, -26186, -24068, -20395, -18195, -11552, -7394, -4623, 
    200, 3362, 9808, 12568, 17445, 19957, 22737, 26311, 28388, 30085, 30068, 
    30304, 31585, 29665, 28837, 27014, 24622, 19480, 15892, 11249, 9674, 
    4543, -473, -3003, -8181, -13744, -17437, -21181, -23899, -25233, -28416, 
    -29917, -30318, -32299, -29817, -29113, -27901, -26521, -23917, -21137, 
    -18685, -13616, -9668, -5380, -1693, 4865, 7546, 14017, 16495, 21038, 
    23912, 24499, 26808, 29553, 31344, 32170, 30004, 30003, 28436, 25829, 
    24698, 20468, 16565, 13545, 9568, 5182, 395, -4425, -8114, -12824, 
    -14940, -19323, -24642, -24696, -27713, -29574, -31389, -30692, -30326, 
    -29644, -27989, -26139, -23394, -20135, -17747, -14230, -9955, -5775, 
    -655, 3030, 8820, 10922, 14564, 20624, 22680, 24526, 27662, 30134, 30249, 
    30940, 30517, 30447, 29107, 26907, 22888, 21792, 18228, 14047, 11236, 
    6141, 939, -2413, -7499, -11868, -17398, -20186, -22580, -25159, -26932, 
    -27885, -29652, -30937, -28832, -30345, -29834, -25853, -23638, -21315, 
    -18849, -14473, -8902, -6262, -2899, 4128, 6143, 10266, 15037, 19029, 
    23129, 25835, 27600, 28947, 30258, 31215, 30537, 30098, 27838, 25979, 
    23394, 22412, 17652, 13319, 10808, 6561, 2520, -2677, -5455, -12676, 
    -15503, -19157, -22093, -26149, -26353, -29761, -28708, -30439, -30873, 
    -30026, -27807, -28401, -24807, -20714, -17625, -15792, -11528, -4888, 
    -1718, 3460, 7074, 11594, 15494, 17862, 20576, 25616, 27427, 28391, 
    28966, 30351, 31366, 29066, 29808, 27455, 25790, 21446, 17837, 14621, 
    10203, 6343, 573, -1080, -6739, -10371, -14630, -18435, -21783, -24768, 
    -26864, -29081, -29075, -30885, -29009, -30206, -28023, -26620, -26240, 
    -21586, -17334, -15450, -11368, -6076, -2175, 2080, 5866, 10352, 14605, 
    17791, 20335, 24620, 27797, 30522, 29589, 30584, 30507, 29168, 27342, 
    27835, 25585, 21278, 17171, 15605, 12380, 7779, 1444, -1172, -6589, 
    -10686, -13634, -18807, -22174, -22799, -27705, -29142, -29560, -31242, 
    -31169, -29816, -29813, -27035, -25166, -22787, -19566, -16038, -12004, 
    -6590, -3558, 1663, 7108, 10485, 14625, 19717, 21038, 24660, 28328, 
    28983, 28642, 31187, 30959, 30230, 28878, 27823, 24021, 22400, 19456, 
    15073, 12152, 7016, 3775, -1118, -7181, -8876, -15201, -17766, -20295, 
    -24558, -26621, -28620, -29132, -30967, -31178, -30098, -29027, -27314, 
    -23681, -23193, -19291, -16036, -12180, -9184, -3642, 793, 6132, 11271, 
    13701, 17668, 20785, 23719, 26210, 27670, 30350, 29898, 30611, 29806, 
    29176, 28383, 23767, 23635, 20146, 15355, 11827, 8340, 2686, -550, -5405, 
    -7984, -13405, -17791, -20289, -25522, -26366, -27440, -29280, -29794, 
    -30304, -30282, -29644, -27253, -24528, -22725, -19867, -16439, -12770, 
    -7585, -3506, 517, 5841, 11164, 13232, 18458, 20861, 24167, 25998, 27806, 
    29478, 31613, 30576, 30173, 29554, 28279, 26092, 21828, 19287, 16438, 
    13021, 6886, 5176, -121, -4438, -8441, -12813, -17680, -21192, -24764, 
    -26101, -29256, -29071, -31928, -30135, -29577, -30563, -26633, -25450, 
    -23840, -19340, -16173, -10623, -8886, -5009, -316, 3906, 9199, 13094, 
    16110, 21199, 24928, 25613, 28141, 28657, 31344, 31380, 29291, 30431, 
    26927, 25583, 22731, 20390, 15433, 11877, 7776, 4191, 386, -4454, -9804, 
    -13106, -17910, -20745, -22328, -26931, -26912, -28472, -31258, -29831, 
    -29637, -28448, -29393, -25658, -21867, -20584, -15782, -12336, -9784, 
    -4886, -487, 4760, 9814, 12188, 16349, 19235, 22907, 27084, 28548, 27999, 
    31651, 30610, 30732, 29213, 28747, 25780, 24213, 19078, 17220, 13218, 
    7862, 4702, 1537, -5454, -9122, -11669, -16814, -19694, -22919, -26218, 
    -29221, -30236, -30116, -31641, -29758, -30761, -28853, -26983, -23027, 
    -20526, -15787, -13542, -10232, -2939, -101, 3877, 9681, 12421, 15929, 
    18010, 23623, 25469, 29254, 29812, 30458, 31735, 31718, 29369, 29485, 
    27100, 24213, 20424, 17394, 13150, 8065, 4591, 1279, -2811, -7514, 
    -12510, -14991, -18786, -24529, -26024, -27966, -28627, -29362, -31345, 
    -30318, -28494, -28418, -25773, -24073, -21253, -17440, -13628, -10088, 
    -4866, -867, 2655, 7379, 12448, 14460, 20169, 22221, 26407, 27633, 29184, 
    29756, 29111, 30127, 29563, 27361, 25937, 24347, 20790, 17769, 12248, 
    9687, 4195, 1212, -2754, -7563, -10406, -14382, -20168, -23099, -26460, 
    -27579, -29767, -30606, -30573, -30883, -29604, -27772, -26670, -23511, 
    -22158, -18177, -13496, -10119, -6157, -1048, 3413, 6748, 12619, 16082, 
    19526, 22857, 26289, 26173, 29373, 30208, 31399, 31008, 29808, 29823, 
    26894, 23306, 20302, 18075, 14659, 10240, 5652, 2652, -1396, -7275, 
    -12415, -15891, -19522, -21552, -23450, -26733, -29689, -29224, -30164, 
    -30735, -28819, -28993, -27714, -25530, -22300, -17234, -13772, -9631, 
    -7569, -602, 3855, 6160, 11651, 15087, 19375, 22623, 24952, 26367, 29481, 
    31097, 30038, 31219, 29358, 28712, 27307, 23362, 21230, 18823, 15059, 
    10431, 7881, 2223, -1173, -6207, -11355, -15534, -18151, -21825, -26359, 
    -25670, -29816, -31155, -29854, -29892, -30396, -29559, -25367, -24991, 
    -21284, -17881, -13522, -10395, -5811, -2935, 2756, 6725, 10582, 14086, 
    19192, 22188, 24304, 25984, 29165, 29813, 29459, 30818, 29937, 27442, 
    28489, 24740, 21982, 19807, 16220, 10980, 6901, 2490, -2517, -6235, 
    -10241, -14696, -18028, -21264, -25627, -26252, -29583, -29385, -30382, 
    -30608, -30559, -29438, -27805, -25926, -20663, -20434, -15278, -11346, 
    -8049, -3527, 1236, 6420, 10433, 14490, 18359, 20403, 24512, 25592, 
    28937, 30534, 30149, 32271, 30719, 30733, 27074, 25326, 22282, 20050, 
    15007, 12797, 7320, 4635, -1822, -6990, -10322, -15311, -19303, -21180, 
    -23050, -26647, -29296, -29502, -32206, -29651, -31502, -28944, -27862, 
    -25563, -21906, -19611, -14999, -11549, -6082, -2365, 1629, 5387, 9355, 
    14283, 17457, 20094, 23593, 26805, 28069, 29132, 30673, 31429, 28637, 
    28061, 27228, 25728, 22038, 19229, 15066, 12822, 8078, 2571, -1587, 
    -5654, -9287, -13597, -18276, -20331, -25638, -26255, -29548, -29090, 
    -30796, -30487, -30636, -29025, -27018, -26018, -22922, -19901, -15839, 
    -11703, -7353, -3258, 1969, 4917, 9031, 13071, 17127, 19759, 22350, 
    26174, 27810, 30606, 29201, 29381, 29893, 29071, 29070, 24128, 23599, 
    20530, 17690, 11010, 9088, 1858, -1587, -5024, -7764, -13709, -17534, 
    -20555, -22457, -25247, -27278, -30653, -29939, -30699, -29739, -28158, 
    -26818, -25122, -24790, -20287, -17151, -12232, -8158, -3933, -285, 5944, 
    8913, 12778, 16441, 20309, 22983, 26058, 28324, 29132, 30400, 30228, 
    31797, 30495, 28257, 24241, 21871, 19442, 17987, 12977, 9611, 3119, -259, 
    -4577, -8509, -12708, -17116, -21230, -24145, -26573, -27822, -29748, 
    -30234, -29317, -30990, -29434, -28553, -25202, -23421, -20861, -15611, 
    -13831, -10084, -4079, 802, 5115, 9705, 11992, 16622, 19697, 23343, 
    25602, 28991, 30350, 30435, 30583, 31354, 29231, 28701, 27279, 23101, 
    19249, 18092, 12682, 8076, 4442, -447, -3663, -8310, -11313, -15906, 
    -20045, -23247, -26758, -28337, -28896, -29741, -30754, -31559, -30635, 
    -29529, -24878, -23084, -20200, -18519, -12644, -7794, -6143, -911, 3978, 
    8579, 11531, 16517, 20633, 22348, 24819, 28247, 30438, 30651, 29975, 
    31417, 31035, 29517, 25316, 24297, 20782, 16547, 13539, 9219, 5219, -99, 
    -3249, -7879, -11505, -17384, -18153, -23050, -24710, -28882, -28615, 
    -29022, -29788, -30322, -28428, -27627, -26864, -23221, -20989, -18682, 
    -13427, -10320, -6848, -1971, 2123, 7511, 11705, 15322, 18396, 22976, 
    24299, 26822, 29674, 31340, 31048, 30790, 31528, 28991, 25317, 23274, 
    21407, 16630, 14025, 11270, 5605, 997, -4280, -8609, -10749, -16427, 
    -19968, -22190, -25149, -28464, -28705, -30801, -30071, -31190, -28844, 
    -28255, -26864, -25162, -20598, -18407, -14058, -10382, -4796, -1134, 
    1527, 7525, 11065, 14867, 19251, 21167, 26379, 26600, 29942, 28898, 
    31500, 29423, 29757, 30004, 25992, 24317, 21291, 18673, 14197, 10170, 
    5504, 1787, -2612, -5948, -12241, -15762, -17905, -21146, -25064, -27395, 
    -29971, -30436, -30077, -31377, -31045, -28491, -26227, -23793, -21577, 
    -17024, -13821, -10553, -6567, -1973, 2608, 6340, 10494, 15549, 19517, 
    23381, 26111, 27039, 27906, 29983, 31075, 29196, 29609, 29406, 27255, 
    23909, 21416, 19635, 15894, 11052, 5014, 1968, -1928, -6561, -10371, 
    -15676, -20372, -21434, -23956, -26235, -28699, -30163, -30934, -29573, 
    -31024, -28905, -27633, -24974, -21248, -18342, -14444, -11026, -8066, 
    -2354, 1749, 7189, 10959, 15679, 17170, 22882, 25065, 26965, 29040, 
    30229, 30315, 30374, 29069, 30256, 27468, 25161, 21105, 18047, 16606, 
    12051, 6323, 1571, -1892, -7130, -9728, -15893, -18033, -21392, -24850, 
    -27183, -29079, -30513, -29176, -30742, -29662, -28384, -27361, -24569, 
    -23169, -19165, -13820, -11494, -7448, -1894, 1959, 5784, 8860, 14243, 
    19097, 22151, 23257, 25854, 28160, 31312, 30746, 31419, 30387, 30219, 
    28045, 24509, 20883, 18456, 14547, 10934, 5398, 2019, -371, -6663, -9596, 
    -14030, -16669, -22191, -26093, -28164, -28930, -30007, -31365, -31942, 
    -31553, -29160, -27474, -24894, -23828, -19648, -15762, -11546, -6854, 
    -4068, 1630, 5930, 10321, 15089, 18695, 21791, 24213, 26576, 28312, 
    30345, 30708, 32234, 30309, 28948, 27801, 25158, 22928, 19847, 15153, 
    13195, 8472, 2792, -1988, -3741, -10307, -14285, -16063, -20708, -23324, 
    -27127, -27260, -29201, -30320, -31971, -30724, -28710, -29080, -24427, 
    -23126, -18619, -16946, -11582, -6880, -3257, 334, 5523, 9995, 13168, 
    15747, 22554, 23996, 26005, 28109, 30154, 30406, 31084, 31206, 29117, 
    28495, 24777, 21309, 19106, 15742, 12450, 7204, 3459, 52, -5923, -10380, 
    -13249, -16636, -20371, -23634, -26830, -28460, -29395, -30449, -31781, 
    -29874, -29654, -27987, -25513, -21748, -21016, -15692, -12228, -9287, 
    -3384, 238, 3415, 10229, 13319, 16375, 21024, 24997, 26512, 27989, 29643, 
    30660, 30737, 30341, 31162, 28230, 26001, 22817, 21803, 16884, 13113, 
    9740, 3252, -1105, -4645, -8018, -13449, -16789, -21149, -23240, -24561, 
    -27510, -27949, -30764, -31482, -28994, -30676, -28366, -27003, -22916, 
    -20589, -17351, -14278, -8547, -3977, -751, 3867, 8613, 13565, 16963, 
    20408, 23991, 27524, 28240, 29199, 31151, 30533, 30033, 29459, 27969, 
    25112, 24588, 21361, 15788, 11753, 9077, 6011, 956, -5027, -8938, -12090, 
    -16615, -19693, -24547, -25663, -28752, -29617, -29803, -31725, -31976, 
    -29611, -27721, -27092, -22959, -19957, -16873, -13269, -9136, -4246, 
    -772, 4973, 6443, 11286, 16747, 19417, 23025, 26352, 26505, 29815, 30128, 
    31549, 29824, 29421, 27836, 25459, 24248, 20518, 16716, 12974, 9267, 
    5197, -104, -3686, -9393, -11668, -16231, -19721, -22589, -26459, -28186, 
    -29221, -31015, -29745, -30384, -28960, -27636, -24690, -23745, -22060, 
    -18756, -13969, -10276, -5654, -1827, 4065, 6978, 12748, 16300, 18182, 
    24267, 26266, 26508, 29755, 31425, 31583, 31787, 31041, 28777, 27096, 
    23762, 21198, 17567, 13697, 8350, 5348, 598, -2025, -6931, -11650, 
    -16560, -19545, -23050, -24852, -27365, -27863, -31141, -31417, -30462, 
    -30226, -27501, -27139, -24223, -22038, -18643, -14292, -10593, -5295, 
    -593, 2661, 7372, 13025, 15561, 19778, 22431, 24676, 28755, 28517, 29576, 
    29355, 29797, 31403, 27902, 27578, 25015, 19721, 17368, 14162, 9985, 
    6111, 1892, -2515, -7704, -10314, -14762, -19529, -21899, -23668, -26405, 
    -30166, -30468, -30789, -32041, -30672, -28440, -25338, -24118, -21028, 
    -18421, -12975, -11329, -5300, -3042, 3130, 7624, 10417, 15230, 19631, 
    21982, 24129, 28556, 28363, 29459, 30175, 31327, 30587, 28876, 26184, 
    24903, 20987, 19378, 14848, 9301, 7189, 2099, -3514, -7095, -11011, 
    -13741, -20317, -22449, -24740, -27174, -28414, -29958, -30891, -31268, 
    -30304, -29960, -25749, -24217, -22907, -16551, -13877, -10301, -5210, 
    -2629, 2946, 7363, 10633, 15758, 17712, 22755, 25357, 27145, 27604, 
    30459, 31683, 30227, 29315, 30468, 27620, 25492, 21040, 18178, 14853, 
    11327, 6953, 2127, -2348, -5789, -11391, -14677, -19589, -19846, -23485, 
    -27280, -29919, -28863, -30054, -31575, -31540, -29023, -26510, -25196, 
    -23785, -18323, -15230, -9976, -6533, -3660, 107, 6059, 11100, 13908, 
    18640, 20637, 23696, 26795, 28927, 31519, 32427, 31428, 30002, 28190, 
    27771, 24259, 22217, 19294, 15612, 11980, 6403, 4232, -2763, -4969, 
    -10619, -15844, -17100, -21044, -25353, -26177, -28537, -28656, -30105, 
    -31818, -29668, -29321, -27067, -24998, -21400, -19366, -14885, -10462, 
    -6103, -2377, 1, 6612, 10014, 12408, 17649, 21372, 22524, 27346, 27813, 
    29886, 30237, 30508, 31484, 29089, 26158, 27163, 22537, 19481, 14409, 
    13594, 6824, 4428, -1503, -5863, -9296, -13873, -16286, -22496, -25825, 
    -25947, -27167, -29677, -29463, -32403, -30978, -27723, -28599, -24466, 
    -23057, -18834, -16086, -10780, -9366, -3533, 436, 4863, 9086, 13606, 
    17195, 20840, 24845, 26178, 29613, 31019, 31779, 31608, 31039, 31037, 
    28213, 26244, 22087, 19543, 16851, 12694, 6934, 3860, -612, -3969, -9873, 
    -13281, -16679, -21367, -23952, -26721, -29673, -30212, -30386, -30226, 
    -30596, -28408, -27131, -25686, -22959, -21374, -16207, -12536, -7220, 
    -4410, 1428, 3881, 8042, 14566, 15849, 19817, 24357, 25452, 29227, 30817, 
    30521, 31864, 31746, 30709, 27607, 25339, 23095, 19200, 17740, 12621, 
    9284, 4145, -790, -5133, -7818, -13142, -16485, -19488, -22750, -26498, 
    -29379, -29927, -31089, -29656, -29647, -30277, -26578, -26929, -22785, 
    -20184, -17369, -12447, -7773, -4560, 903, 4446, 10278, 13318, 16148, 
    20791, 23283, 25247, 29151, 30384, 30864, 30563, 29939, 29124, 26988, 
    26423, 23704, 19216, 18410, 14216, 8674, 4173, -1097, -5183, -8565, 
    -13698, -17621, -19976, -22333, -25299, -27222, -27992, -30066, -30667, 
    -31528, -28449, -28947, -25863, -23586, -21336, -16167, -12842, -10265, 
    -4420, -375, 4760, 6660, 12731, 16423, 18426, 22472, 25963, 27889, 30890, 
    30963, 30090, 31305, 28932, 27118, 27139, 24833, 21118, 18293, 13859, 
    9230, 4180, 904, -5040, -7985, -11791, -15674, -18548, -21297, -25964, 
    -27060, -29410, -28914, -31079, -30918, -29872, -26986, -25173, -24026, 
    -20028, -17182, -13181, -8641, -6305, -175, 3550, 7428, 12177, 15710, 
    18717, 22697, 24377, 27326, 29875, 30337, 30526, 29589, 31194, 29129, 
    27557, 22974, 22531, 17669, 12649, 9904, 5475, 2645, -2988, -6412, 
    -12324, -15613, -20568, -22458, -25670, -27562, -28576, -29827, -31217, 
    -30450, -28578, -28389, -27031, -24905, -20056, -17861, -13767, -9207, 
    -6212, -2499, 2712, 7528, 10419, 14338, 18773, 21569, 24777, 27938, 
    28741, 31161, 31559, 31450, 29772, 28546, 26712, 23878, 19803, 17987, 
    13432, 10873, 5761, 1253, -2985, -7587, -11057, -14961, -19715, -21620, 
    -25476, -26293, -28251, -29703, -31277, -30676, -30015, -29973, -26093, 
    -22540, -22683, -17181, -16019, -9908, -7460, -2450, 1661, 7827, 11884, 
    13984, 19175, 21635, 26282, 27412, 28080, 29354, 31937, 30291, 30457, 
    28210, 28413, 24637, 21819, 17805, 15426, 9715, 5663, 1644, -2070, -6443, 
    -10927, -16585, -19898, -20123, -24766, -28111, -27956, -30258, -31142, 
    -32187, -29245, -29266, -28244, -25916, -21835, -18963, -13537, -11176, 
    -5674, -2668, 2882, 6683, 11053, 15332, 18328, 22428, 25226, 28494, 
    28367, 28496, 30406, 30153, 30766, 27452, 27086, 24464, 22485, 17972, 
    16105, 10732, 6975, 2744, -1583, -6514, -11654, -12830, -18764, -22337, 
    -23966, -26893, -28382, -29212, -30657, -30427, -30412, -28798, -27091, 
    -25778, -23083, -18213, -14741, -9793, -5354, -3060, 3388, 6579, 11378, 
    13289, 18009, 21763, 24833, 26928, 28216, 29953, 30034, 30236, 30348, 
    30157, 28150, 25248, 21347, 18549, 14571, 12382, 6542, 2679, -1379, 
    -6748, -9544, -14844, -17003, -21979, -23871, -26574, -28535, -29439, 
    -30417, -30435, -31730, -29230, -27557, -26371, -22327, -19001, -15457, 
    -10705, -7776, -2655, 1215, 6675, 8716, 13084, 16765, 20435, 24955, 
    28037, 27964, 30270, 30387, 32271, 31173, 29073, 27070, 25802, 22321, 
    19119, 14405, 11731, 7149, 1511, -373, -6278, -9430, -14352, -18364, 
    -20026, -23497, -25791, -27218, -31127, -31067, -30986, -30385, -28782, 
    -29184, -25200, -21856, -19829, -16706, -12139, -9086, -3915, -477, 4579, 
    9253, 14810, 16424, 20583, 23025, 25917, 28914, 29757, 30888, 29894, 
    29473, 30411, 28747, 25341, 22239, 18627, 16348, 12304, 8481, 3511, 518, 
    -5817, -9903, -13962, -16609, -19769, -22306, -26278, -28931, -30230, 
    -29235, -30581, -29876, -29002, -29319, -26315, -23606, -18879, -17707, 
    -12566, -8610, -3907, 468, 5411, 8090, 13010, 16462, 19698, 24183, 24886, 
    28176, 28923, 31747, 30596, 30519, 29382, 27553, 24516, 22211, 20556, 
    18246, 12014, 7333, 3373, -1192, -3688, -8459, -13225, -17886, -20423, 
    -22944, -26271, -28831, -29092, -31412, -31989, -30329, -31280, -28758, 
    -26877, -24824, -21733, -17116, -12327, -9868, -5393, 551, 3174, 8134, 
    11318, 15653, 21628, 21820, 27411, 28586, 30242, 30511, 30539, 31803, 
    29961, 27701, 26006, 22973, 20126, 16470, 13925, 8962, 5012, 99, -4005, 
    -7137, -12699, -16981, -20946, -22764, -25978, -27372, -30056, -31412, 
    -29790, -30987, -29961, -28142, -25584, -23950, -20388, -16747, -13799, 
    -8481, -5112, 1005, 4397, 7437, 11382, 15195, 19900, 22300, 25453, 28698, 
    27790, 31729, 29674, 31023, 29166, 30065, 26789, 23618, 20163, 16550, 
    13210, 10787, 4870, 96, -3971, -6966, -12653, -16795, -20436, -21412, 
    -25834, -27915, -29544, -29121, -31417, -29276, -31239, -28732, -27689, 
    -23092, -21370, -17943, -14272, -9701, -3893, -1717, 4642, 7390, 12914, 
    15490, 19407, 22565, 26271, 27848, 29438, 30889, 30862, 29668, 30006, 
    28252, 27466, 23747, 21211, 18082, 14724, 10829, 5839, 1037, -4975, 
    -6809, -12273, -15267, -20980, -21114, -25188, -27049, -28204, -30296, 
    -30130, -30081, -29745, -29784, -25262, -23202, -19894, -16544, -14878, 
    -9504, -5610, -686, 3405, 8809, 11357, 14413, 18753, 22241, 23366, 28768, 
    29936, 30875, 30717, 32257, 30633, 27522, 25525, 23171, 20881, 18554, 
    15094, 9863, 7374, 502, -2798, -6556, -13213, -14170, -19311, -23565, 
    -25407, -28740, -27902, -31313, -30925, -30246, -30336, -28356, -26496, 
    -25598, -23136, -17737, -14410, -9227, -6908, -643, 2967, 5561, 10588, 
    16725, 17380, 21646, 25213, 26129, 28259, 28809, 29392, 29513, 28543, 
    30137, 27577, 23085, 22433, 16707, 15428, 11120, 4845, 3012, -3571, 
    -6931, -10058, -14787, -18405, -21468, -25651, -25900, -29224, -29653, 
    -32244, -30771, -29561, -27357, -27209, -24214, -21455, -18367, -13405, 
    -11220, -6839, -1772, 2891, 6874, 9864, 15824, 18301, 21260, 23270, 
    27634, 28895, 29620, 30175, 31625, 30126, 28055, 26099, 24810, 23430, 
    19299, 16056, 9808, 5892, 2020, -1348, -5891, -10410, -15999, -18160, 
    -21659, -24994, -27172, -29460, -29056, -31481, -30044, -30645, -28563, 
    -27541, -25585, -22358, -18907, -14785, -11133, -7274, -1455, 1805, 6677, 
    11690, 13852, 18724, 22643, 23636, 27977, 29038, 29948, 30818, 31006, 
    28637, 28131, 28179, 26093, 21395, 18208, 14654, 11271, 5470, 2204, 
    -2807, -5241, -10756, -14830, -18242, -22077, -25017, -25856, -28839, 
    -29590, -30984, -31187, -29803, -28034, -27731, -24590, -22718, -18366, 
    -15278, -12048, -7966, -2316, 2556, 4939, 9737, 12179, 17633, 21117, 
    23812, 27011, 28627, 28799, 31867, 30690, 30266, 28275, 29358, 24721, 
    22897, 19559, 15551, 11763, 7064, 4368, -1920, -4101, -9757, -13292, 
    -17523, -20314, -23172, -25732, -27533, -29908, -30932, -30429, -30265, 
    -29530, -26358, -25389, -22301, -19475, -14818, -11889, -5998, -3293, 
    1379, 7136, 9327, 13053, 17103, 21258, 23940, 26066, 28237, 29924, 30919, 
    29458, 31131, 30033, 27790, 25509, 22950, 19850, 17180, 13707, 6491, 
    3444, 212, -4559, -10357, -14056, -17891, -20692, -22189, -26509, -27055, 
    -28000, -30473, -31252, -31504, -29246, -26812, -23979, -24176, -20682, 
    -16713, -12699, -7352, -2838, 1807, 3793, 10501, 13008, 17260, 20815, 
    23972, 25714, 28427, 30114, 29974, 31760, 30717, 29312, 26265, 27378, 
    22843, 18554, 16516, 11307, 8253, 5462, 300, -4176, -8779, -12722, 
    -16887, -18536, -22452, -25343, -26275, -30235, -31293, -31798, -30620, 
    -30198, -28725, -26221, -23955, -20351, -16635, -12914, -7897, -4542, 
    -1038, 5913, 10043, 13242, 16595, 19415, 22288, 26935, 28599, 28386, 
    30662, 31871, 31232, 29937, 27922, 25506, 22191, 20496, 16935, 12621, 
    8354, 3201, -761, -4533, -9264, -13897, -16373, -19889, -24609, -26585, 
    -27681, -29796, -30012, -32207, -30033, -29866, -27640, -25532, -24773, 
    -19470, -17370, -13730, -9829, -5781, 267, 4119, 8841, 12072, 15708, 
    20948, 21598, 25980, 27313, 30794, 30909, 30614, 30624, 29521, 27556, 
    26582, 24115, 20265, 16137, 12540, 7757, 5792, 261, -4716, -8203, -10841, 
    -16138, -18962, -22939, -24837, -28547, -30268, -30490, -30768, -30129, 
    -29727, -28793, -25758, -25557, -20968, -18763, -14277, -9442, -6241, 
    -935, 3097, 7107, 12387, 16621, 19912, 22705, 26214, 27963, 29496, 30855, 
    32150, 30680, 30100, 27750, 26650, 24380, 21106, 16917, 13887, 7821, 
    5622, 741, -3072, -5973, -10290, -15775, -18832, -22512, -23448, -28138, 
    -30886, -29424, -32234, -30147, -29710, -28329, -25692, -23371, -21742, 
    -17911, -13138, -10669, -5309, -1760, 3103, 6876, 11178, 15841, 18373, 
    21663, 26184, 28397, 29916, 30484, 30578, 31034, 28864, 27278, 27340, 
    23386, 20310, 18006, 13030, 11128, 5022, 1014, -3320, -7580, -11116, 
    -15082, -17639, -21876, -26308, -27649, -27780, -29636, -31336, -31506, 
    -28959, -29987, -27357, -24041, -20731, -17572, -14205, -11876, -5756, 
    -1602, 2327, 6264, 11875, 16317, 19128, 22007, 24659, 27546, 28825, 
    30687, 31020, 30442, 29765, 28472, 26357, 24050, 21313, 18028, 14173, 
    10120, 5523, 1063, -1719, -6307, -10695, -14957, -18596, -21477, -24278, 
    -26721, -29338, -30517, -29852, -29961, -31000, -27287, -27320, -24093, 
    -21613, -17589, -13623, -10654, -6251, -844, 746, 6812, 10937, 15627, 
    18350, 21214, 25211, 27700, 28883, 29930, 29414, 31497, 29388, 28555, 
    28842, 25321, 21988, 17048, 14008, 10272, 6359, 2526, -1942, -4788, 
    -11756, -14898, -19095, -20908, -24893, -26279, -29271, -30625, -30799, 
    -29605, -29924, -28968, -27912, -24282, -22423, -18464, -16354, -11019, 
    -7964, -3943, 1545, 6779, 9231, 13086, 17230, 21958, 24749, 26566, 29363, 
    30160, 30691, 31207, 31474, 29912, 27172, 24932, 21880, 17602, 15025, 
    9991, 8310, 2464, -1259, -5439, -10279, -14869, -17809, -22495, -24209, 
    -26024, -28782, -28820, -31213, -30179, -32057, -28537, -27546, -26120, 
    -23127, -19573, -16290, -11691, -6119, -1612, 358, 5581, 9310, 14450, 
    17535, 21499, 22941, 26320, 28035, 30570, 29531, 30561, 29881, 28516, 
    28850, 25547, 23148, 19448, 15029, 11148, 7328, 2179, -564, -5289, 
    -11081, -13765, -16421, -21723, -23859, -26311, -28097, -29786, -30923, 
    -30373, -29528, -30687, -27091, -24994, -22012, -19830, -15744, -10378, 
    -7275, -4037, 1278, 5815, 10264, 12791, 16722, 20023, 23397, 26646, 
    28424, 30580, 29510, 31921, 29903, 29059, 27540, 24881, 21274, 19621, 
    15586, 11614, 9085, 3889, -1243, -4892, -8924, -12253, -16047, -19564, 
    -23330, -26606, -28219, -30585, -30179, -31662, -30682, -27638, -26993, 
    -25149, -24245, -20759, -16264, -12451, -8245, -4596, 1250, 5070, 9869, 
    13605, 16134, 20706, 24619, 27004, 29065, 30408, 30675, 30124, 30252, 
    28510, 28059, 24759, 24462, 19813, 16402, 12876, 8022, 4973, -613, -6070, 
    -8958, -14153, -17988, -19724, -24374, -26389, -29258, -29086, -31632, 
    -30922, -30727, -30424, -28791, -26016, -23693, -20346, -15753, -12890, 
    -8523, -4319, 1219, 4751, 8174, 12763, 15142, 21536, 24099, 26450, 27835, 
    29197, 32158, 30283, 29823, 30279, 28104, 26094, 23946, 19645, 16963, 
    13545, 8686, 5336, 500, -4292, -8797, -12756, -17236, -20556, -24258, 
    -26523, -27342, -28991, -29211, -31059, -31461, -28702, -29311, -24565, 
    -24108, -20991, -17762, -13704, -7666, -5750, -747, 4815, 8678, 12886, 
    16437, 20253, 21909, 26882, 27737, 30440, 30438, 30122, 30067, 28753, 
    26707, 25315, 24069, 19157, 17724, 14052, 9653, 4568, -571, -2946, -6329, 
    -12615, -17810, -21048, -23093, -25308, -27523, -29795, -30518, -30719, 
    -30383, -30781, -27047, -25902, -23867, -20425, -17914, -12666, -8981, 
    -5323, -1218, 3832, 9298, 11986, 17227, 20735, 23817, 24119, 26653, 
    29423, 28765, 30997, 31058, 30248, 28324, 27812, 23302, 20849, 18827, 
    13080, 10281, 6398, 586, -2805, -8033, -11010, -15560, -19540, -23881, 
    -24711, -28024, -30850, -29171, -30042, -31672, -30271, -29003, -27186, 
    -24513, -20640, -18052, -13950, -10092, -5688, -1178, 2489, 8385, 11078, 
    15532, 19463, 22531, 25715, 27982, 27383, 30563, 30920, 30975, 30753, 
    28938, 27835, 25843, 21479, 18376, 13233, 9206, 5159, 621, -1725, -8604, 
    -10973, -14492, -20690, -21386, -25429, -26380, -30063, -30128, -31083, 
    -30438, -29545, -28869, -27244, -24257, -21733, -17536, -13937, -9551, 
    -7128, -715, 2662, 8338, 9650, 15946, 18737, 23175, 25527, 27481, 27707, 
    28436, 30709, 30899, 30092, 28891, 26808, 25542, 20903, 17960, 14534, 
    10131, 6756, 2206, -2563, -8021, -9576, -14416, -19608, -20642, -24396, 
    -27969, -28931, -30773, -30920, -30507, -30700, -30397, -27001, -23591, 
    -22064, -18631, -14765, -10036, -7241, -1989, 2170, 7043, 10337, 13571, 
    17981, 21602, 24442, 26821, 29689, 29653, 31881, 31376, 30039, 29685, 
    27797, 24326, 20671, 18005, 15252, 9638, 6402, 2095, -244, -7691, -11924, 
    -14642, -19515, -20963, -24410, -25903, -28323, -29713, -30823, -31590, 
    -30848, -28489, -28423, -25591, -22811, -18781, -15015, -10382, -6938, 
    -1024, 2621, 4389, 9531, 14375, 18211, 21124, 23400, 25287, 27630, 28634, 
    30163, 30422, 30049, 28339, 27591, 24854, 22179, 18451, 14154, 11698, 
    6661, 3953, -2324, -5155, -8749, -14260, -16849, -21826, -24839, -26085, 
    -28666, -28274, -30338, -32487, -31530, -29657, -28121, -26975, -21328, 
    -18909, -16431, -9755, -7208, -3285, 1219, 4422, 10823, 14251, 16265, 
    21533, 23720, 26527, 26950, 29502, 31848, 30777, 30232, 30713, 27689, 
    26595, 22361, 18953, 14222, 12592, 5858, 3493, 471, -6769, -10807, 
    -12929, -15999, -19506, -24446, -26137, -28633, -28614, -29639, -30881, 
    -31093, -28254, -27002, -25177, -22488, -20558, -15590, -12325, -8314, 
    -2846, 1537, 5320, 8797, 12577, 18015, 21248, 23049, 27339, 28722, 29274, 
    30790, 29153, 29967, 29349, 27346, 25290, 22517, 20529, 16178, 12503, 
    9352, 4211, -892, -3937, -9957, -14066, -17344, -19759, -24727, -25869, 
    -28243, -30359, -30440, -31415, -29241, -29847, -26789, -25947, -23297, 
    -19610, -15494, -12955, -7531, -2836, 473, 4459, 9272, 13636, 18018, 
    20891, 24414, 27335, 27305, 29730, 31561, 30294, 29935, 29429, 27770, 
    25536, 23035, 20908, 17333, 13055, 9185, 5450, 567, -4257, -8699, -13000, 
    -17401, -19890, -24000, -26617, -28528, -29679, -31518, -30906, -30118, 
    -28425, -27030, -26125, -23272, -19937, -16241, -12568, -9025, -5278, 
    -10, 4926, 8233, 11977, 17579, 18656, 21492, 26468, 28898, 29327, 31312, 
    31376, 31705, 29525, 28077, 25696, 23481, 19097, 17750, 14348, 7965, 
    5504, -507, -2899, -7493, -12792, -17260, -18521, -23639, -25204, -27825, 
    -28569, -30614, -29332, -30315, -30733, -28412, -26096, -23631, -20338, 
    -15953, -12609, -8968, -5319, -1078, 4057, 9174, 12310, 17060, 18741, 
    22246, 25968, 26826, 28280, 30274, 31189, 31000, 29097, 26568, 25604, 
    24118, 19460, 18129, 13448, 9245, 6195, -93, -3051, -8056, -13365, 
    -15949, -19997, -23151, -25892, -28255, -29052, -30646, -31574, -30716, 
    -28629, -28819, -27149, -23092, -21373, -17951, -13863, -8330, -5337, 
    -2085, 4803, 6877, 11953, 15447, 19898, 23486, 24879, 26886, 29236, 
    30165, 31070, 31871, 29653, 29320, 26046, 25018, 19775, 19144, 14072, 
    9313, 5290, 1415, -1882, -7477, -10820, -15950, -19869, -21549, -25602, 
    -29080, -27897, -28956, -30206, -31306, -30230, -27610, -27407, -23865, 
    -21044, -19048, -15780, -8676, -4328, -7, 3305, 7669, 11970, 15315, 
    19026, 21887, 25862, 27501, 29690, 30110, 31457, 31226, 29606, 29123, 
    25800, 24686, 22115, 18378, 14389, 9922, 5929, 2458, -2250, -6390, 
    -10825, -15581, -19989, -21170, -24906, -28339, -29288, -28411, -31549, 
    -30376, -29329, -30417, -25979, -22590, -20672, -17723, -14325, -10390, 
    -5226, -1032, 3168, 6405, 12270, 15587, 18180, 20623, 24926, 26599, 
    29475, 29885, 29892, 30070, 30298, 28632, 27905, 24006, 21882, 18403, 
    13769, 11063, 8084, 3047, -3504, -7927, -11435, -13543, -18850, -22246, 
    -23930, -26900, -28829, -31491, -31657, -30025, -29757, -29134, -25705, 
    -25083, -21533, -16952, -15885, -11380, -7169, -1532, 2068, 7689, 10090, 
    15518, 17463, 21905, 24035, 26058, 29998, 30726, 30217, 30681, 29887, 
    30002, 27949, 25850, 21593, 18844, 15182, 11051, 7296, 1204, -572, -5497, 
    -11619, -13949, -17938, -21859, -24588, -25220, -29154, -30984, -29723, 
    -30506, -29378, -29058, -26628, -24632, -21998, -19775, -16657, -12112, 
    -7986, -2572, 1174, 7725, 11626, 14277, 17183, 20986, 23758, 27900, 
    29077, 29810, 29887, 29387, 30345, 29851, 27155, 26391, 22824, 19606, 
    15426, 11937, 8473, 2514, -1001, -4098, -10603, -14335, -16928, -21163, 
    -23592, -28372, -28784, -30313, -30318, -30877, -31804, -29867, -27731, 
    -25491, -22920, -19485, -15565, -13339, -7147, -3504, 482, 6782, 10112, 
    13934, 17553, 21060, 23236, 26109, 28925, 29806, 30134, 30252, 30362, 
    29308, 27461, 25396, 23501, 19757, 16253, 12791, 8111, 1973, -1689, 
    -5159, -9585, -13604, -19064, -21407, -23413, -28243, -28978, -29379, 
    -32490, -32075, -31373, -28451, -29198, -26043, -23788, -19492, -16012, 
    -10443, -7278, -3848, 1455, 5633, 10076, 14197, 17933, 20465, 23531, 
    25157, 28076, 30450, 30084, 31052, 29437, 29963, 28086, 26297, 22456, 
    19755, 15590, 12198, 7131, 2289, 871, -5508, -10106, -14632, -15664, 
    -20462, -24330, -27010, -27469, -30308, -31051, -30775, -29724, -28074, 
    -27322, -23820, -21321, -20592, -16454, -13523, -8364, -3694, -568, 3432, 
    10282, 14436, 17490, 20761, 22720, 26980, 28394, 29358, 30124, 30172, 
    29526, 29309, 27417, 26056, 21575, 19371, 17683, 12230, 7667, 4480, -144, 
    -4576, -8977, -13735, -15807, -19556, -24695, -26146, -28212, -30085, 
    -29949, -31219, -29512, -28581, -29404, -26850, -24088, -20431, -16993, 
    -11601, -8284, -4594, -1102, 4849, 9521, 13253, 17354, 18805, 22171, 
    25201, 27979, 30098, 30872, 31036, 30389, 29331, 28323, 25950, 23570, 
    20907, 15570, 12196, 7433, 5769, -73, -4332, -7324, -12008, -16239, 
    -18814, -23670, -25602, -28330, -29235, -30929, -30315, -30577, -30683, 
    -28259, -26615, -22909, -19238, -16772, -13127, -7724, -5129, -901, 3373, 
    9962, 11507, 16447, 19695, 22605, 26129, 27193, 28441, 29739, 30527, 
    30269, 29060, 27403, 26275, 23419, 20280, 17751, 13583, 9164, 4756, 1646, 
    -3844, -8440, -11620, -14554, -19132, -22483, -25444, -26892, -29301, 
    -30395, -30439, -30473, -29098, -29735, -27848, -22012, -20246, -17628, 
    -13094, -9722, -6644, -1389, 3011, 6418, 12834, 14578, 20085, 21632, 
    26450, 26434, 29187, 30596, 30243, 31917, 30216, 29041, 26448, 24608, 
    20958, 18027, 14788, 10106, 4173, 938, -4081, -6416, -10625, -17006, 
    -18698, -22281, -24056, -28361, -28897, -30401, -31345, -31316, -29469, 
    -28214, -26364, -23999, -20864, -18592, -15084, -10009, -5897, -2511, 
    2580, 6224, 10158, 15088, 18217, 22435, 25480, 27295, 29483, 29646, 
    29771, 30651, 30747, 29816, 26520, 23778, 20174, 17312, 13133, 10485, 
    7305, 1666, -3454, -8297, -11873, -13776, -17772, -22478, -26602, -27096, 
    -29940, -30679, -30325, -29624, -30793, -29257, -26222, -23099, -21843, 
    -18583, -14899, -11137, -5673, -3025, 2819, 5870, 10524, 13372, 19597, 
    22560, 25217, 27427, 28848, 29937, 31127, 31057, 29498, 29617, 26295, 
    24036, 21890, 19701, 14174, 9816, 8112, 2493, -1629, -6180, -9096, 
    -14971, -18133, -21532, -24747, -27315, -28831, -30864, -30648, -31911, 
    -29731, -29955, -28232, -24159, -21354, -17664, -13861, -11839, -6435, 
    -1279, 1367, 7953, 10876, 14095, 18832, 21647, 24119, 26558, 29028, 
    30165, 31067, 32149, 30441, 28701, 27827, 24472, 22049, 18337, 15260, 
    12450, 6133, 2642, -1880, -6178, -10389, -15202, -19101, -20145, -25521, 
    -26631, -29493, -29334, -31022, -29956, -29267, -28957, -26726, -25200, 
    -21242, -18808, -15084, -10474, -6264, -2306, 861, 6565, 10303, 14858, 
    17943, 20884, 23971, 26218, 27497, 30442, 32335, 29481, 30823, 30057, 
    27727, 24718, 22495, 17714, 15809, 11230, 7272, 3327, -2266, -5385, 
    -9720, -13062, -17968, -21072, -24259, -27245, -29701, -30291, -31122, 
    -30971, -30375, -29171, -28186, -25728, -22088, -18448, -16354, -10902, 
    -7087, -4008, 982, 7165, 10094, 12719, 18900, 20066, 24620, 25060, 29919, 
    29826, 29159, 30434, 30249, 29660, 28407, 25154, 21095, 20515, 17387, 
    11525, 8582, 4782, -904, -6250, -9429, -13606, -18648, -21623, -24697, 
    -26311, -29253, -29969, -31740, -31891, -29998, -29315, -27595, -25790, 
    -22645, -20871, -17102, -11362, -7813, -3287, 1703, 5151, 9444, 14104, 
    17632, 21909, 24052, 25385, 27159, 31134, 31140, 32042, 31478, 29535, 
    27474, 24677, 22740, 19783, 15518, 11973, 9758, 4755, 222, -6181, -10214, 
    -13818, -17520, -20282, -22616, -26157, -26989, -30520, -31570, -31088, 
    -29240, -29546, -28058, -25557, -23645, -20038, -16138, -11308, -7639, 
    -4592, 200, 4769, 8459, 13144, 16963, 20342, 23809, 27509, 28145, 29725, 
    30286, 31406, 29084, 28967, 28004, 25744, 24606, 19784, 16288, 11977, 
    8589, 4305, -1257, -5121, -7394, -11887, -16955, -19901, -23016, -25600, 
    -27998, -29126, -30268, -30841, -30366, -29813, -27831, -25349, -22390, 
    -20762, -15699, -12915, -7935, -5626, -1050, 2546, 8696, 12276, 17724, 
    21365, 22267, 25579, 28121, 28995, 31702, 29773, 30661, 28830, 28906, 
    25360, 24251, 21373, 17465, 12866, 9548, 5312, 709, -3893, -9065, -13082, 
    -16013, -19736, -22791, -25327, -27993, -28992, -30102, -30584, -32353, 
    -28673, -27298, -26183, -23357, -19566, -16293, -13367, -8758, -4928, 
    -285, 3280, 7431, 13209, 17109, 18699, 22967, 26247, 28889, 30134, 31303, 
    30300, 30917, 29601, 28395, 26914, 23322, 20495, 18296, 12751, 10500, 
    5591, 1749, -3027, -8073, -10850, -17157, -19613, -23046, -24059, -29283, 
    -29404, -30267, -30344, -30821, -30396, -28656, -24946, -22085, -21003, 
    -17810, -13130, -9746, -4102, -972, 4438, 6951, 13236, 16285, 19503, 
    23039, 26017, 29412, 29165, 30000, 31458, 31903, 30814, 26980, 26300, 
    24973, 21744, 17153, 14498, 10305, 5143, 721, -2080, -8923, -13104, 
    -15992, -18771, -22454, -26850, -28035, -27986, -29490, -30795, -32044, 
    -29218, -28302, -27571, -24545, -21428, -17274, -15067, -9568, -4700, 
    -1297, 3409, 7830, 10771, 15860, 19044, 22491, 25059, 27585, 29041, 
    29874, 29655, 31674, 30065, 28036, 26683, 23003, 20337, 18412, 15725, 
    10121, 6124, 3193, -3330, -6550, -12619, -16718, -19053, -22781, -24740, 
    -27345, -29237, -31058, -29900, -30519, -30994, -29149, -27694, -24219, 
    -20454, -18736, -14238, -9722, -7555, -1623, 2313, 7553, 12362, 14732, 
    17685, 23337, 24969, 27359, 27942, 29879, 31089, 29949, 29265, 30093, 
    27531, 23548, 22480, 19403, 13849, 10305, 6474, 3073, -2340, -8355, 
    -12354, -15061, -18890, -21259, -25394, -27435, -28300, -28891, -31697, 
    -29793, -28726, -28162, -28570, -24376, -23195, -18353, -13523, -9118, 
    -6730, -2707, 2608, 6422, 10032, 14310, 17893, 22370, 24111, 25940, 
    28459, 28845, 32036, 29418, 30713, 30328, 28686, 25488, 20544, 20221, 
    14546, 10750, 6684, 2587, -2338, -6198, -10423, -14715, -17461, -22922, 
    -25945, -26062, -28258, -31033, -30319, -30718, -29076, -29640, -28542, 
    -23910, -21592, -19167, -16370, -10809, -7316, -2472, 3111, 7135, 10647, 
    14448, 16936, 20953, 26072, 25774, 26865, 29917, 29727, 30688, 28793, 
    27538, 28142, 25618, 22159, 19400, 16412, 12645, 6336, 2649, -1873, 
    -7170, -10848, -13170, -17436, -22293, -25193, -27179, -28764, -29205, 
    -31419, -29919, -28851, -29838, -28369, -25032, -22897, -19087, -14206, 
    -11710, -6765, -2973, 1397, 6132, 10352, 14740, 18469, 20732, 22371, 
    26598, 29096, 30912, 30805, 30683, 30336, 30493, 29045, 25288, 22494, 
    18886, 14545, 12003, 7956, 2448, -452, -6551, -9496, -13303, -18429, 
    -20566, -24612, -24845, -28752, -29104, -29362, -30407, -30837, -29279, 
    -27394, -25911, -24199, -18861, -17093, -12235, -7812, -2300, 559, 5809, 
    9346, 13377, 16481, 20797, 23267, 26737, 27384, 29746, 32094, 32185, 
    29787, 28849, 26763, 24888, 22656, 18728, 15326, 12122, 8700, 4379, -767, 
    -4007, -7741, -12125, -16837, -19936, -24030, -26455, -27704, -28698, 
    -29647, -31303, -29031, -28066, -27955, -25456, -22434, -18822, -14910, 
    -12823, -8556, -2533, -55, 4870, 8686, 13308, 17578, 20172, 23937, 25848, 
    28883, 29371, 31969, 29576, 30545, 29670, 28523, 25621, 22368, 21075, 
    15726, 12245, 9067, 4894, -1703, -4742, -9099, -13339, -15811, -20377, 
    -23611, -25948, -27389, -30053, -30953, -31644, -29331, -29447, -28632, 
    -24689, -22935, -20039, -16743, -12890, -8587, -4542, 917, 3765, 8528, 
    12338, 16170, 19852, 22665, 27185, 29384, 30546, 29580, 31021, 30828, 
    29314, 27863, 26920, 23806, 20026, 17104, 13219, 7487, 4286, 412, -3619, 
    -8594, -13168, -16339, -20759, -22451, -24134, -28276, -30287, -29085, 
    -30802, -29903, -28315, -29633, -26689, -23197, -20105, -16933, -14161, 
    -7809, -5265, 516, 3785, 9791, 12216, 15810, 20443, 22967, 25771, 27355, 
    29990, 29420, 29639, 30426, 29563, 29118, 27239, 23290, 22124, 17146, 
    12959, 8076, 4350, 344, -4758, -7857, -11947, -16550, -20499, -21534, 
    -24250, -28352, -28503, -31103, -31313, -31191, -31311, -28958, -25318, 
    -22398, -21079, -17942, -14749, -9648, -5141, -1804, 1780, 7548, 11635, 
    15036, 19316, 23599, 25232, 27794, 29684, 29868, 30537, 29194, 29897, 
    28662, 26323, 23881, 21646, 16865, 15028, 10361, 5525, 1144, -2770, 
    -7409, -12594, -17350, -19706, -23293, -24099, -28272, -29396, -31075, 
    -30541, -30861, -28798, -28756, -27509, -23635, -22363, -18754, -13467, 
    -11136, -6342, -1778, 3866, 7263, 10464, 16095, 18954, 21659, 25007, 
    28080, 30132, 30672, 30733, 30905, 29049, 28724, 26972, 24154, 22064, 
    19343, 15350, 8284, 5529, 1719, -3318, -7175, -9824, -14940, -17900, 
    -21936, -24255, -29231, -29791, -29075, -30332, -30887, -29527, -28574, 
    -25496, -23032, -21849, -17337, -14597, -9035, -5658, -2036, 3613, 7491, 
    11521, 15648, 17305, 22995, 24543, 26681, 28992, 30223, 29664, 31043, 
    29933, 27367, 26639, 23980, 22022, 18260, 13696, 10066, 5255, 1402, 
    -1427, -5574, -10990, -15187, -19043, -23416, -23106, -27404, -29024, 
    -29282, -31580, -29582, -29710, -28798, -27824, -24607, -23361, -17494, 
    -15680, -12260, -7287, -2926, 2543, 5419, 10182, 16396, 17087, 21020, 
    25077, 27477, 28926, 30142, 31461, 31351, 30485, 27443, 27922, 24004, 
    20281, 17049, 14992, 10955, 6425, 2096, -1079, -6844, -10726, -15455, 
    -17601, -23122, -24078, -26392, -30071, -30795, -31243, -29662, -29226, 
    -28756, -26730, -24528, -21282, -18713, -15208, -10113, -6972, -3528, 
    2911, 5814, 8817, 14888, 17127, 21687, 25098, 26119, 29409, 29631, 29234, 
    30537, 29578, 29495, 27250, 24616, 22100, 18397, 16503, 10184, 6798, 
    2152, -2268, -5547, -10803, -14126, -18163, -20991, -23899, -26819, 
    -29528, -30593, -31500, -31247, -30804, -29198, -28183, -25005, -22593, 
    -20088, -14974, -10944, -7716, -3151, 2, 4215, 9318, 14101, 16794, 21346, 
    25033, 26976, 27782, 31024, 29671, 32012, 30488, 30015, 28298, 24454, 
    23777, 19107, 15933, 11905, 6571, 3371, -2132, -4580, -9348, -12826, 
    -18588, -21553, -24666, -28078, -27475, -28926, -31890, -29226, -31940, 
    -29418, -26064, -25342, -22730, -18918, -15143, -11361, -8780, -3332, 
    -770, 4618, 10997, 14162, 18041, 19076, 23684, 26577, 27586, 29287, 
    30534, 31694, 30288, 28929, 27746, 26194, 21943, 19999, 17086, 12011, 
    8452, 3909, -475, -6487, -10024, -13320, -16984, -20851, -23073, -26671, 
    -28149, -29358, -31681, -30566, -30891, -30707, -27351, -25152, -22765, 
    -19485, -15636, -12528, -8750, -4475, -329, 5585, 7981, 12321, 17195, 
    20777, 21945, 25714, 26978, 28265, 30690, 30601, 30123, 30759, 27729, 
    26288, 22391, 19804, 17558, 13655, 9475, 4302, 80, -3292, -8316, -12938, 
    -17215, -21075, -23471, -26713, -27462, -29585, -30756, -29318, -31218, 
    -30572, -27269, -26090, -21800, -20966, -16042, -11724, -9120, -4918, 
    477, 3354, 9460, 12104, 15741, 19444, 22152, 25502, 28034, 29198, 29951, 
    31396, 29464, 29771, 28401, 25626, 23147, 20219, 15363, 13100, 7876, 
    5251, -748, -5705, -9473, -14091, -17405, -18450, -24173, -25630, -28238, 
    -30226, -29055, -30731, -31254, -29083, -27663, -26326, -23449, -19415, 
    -16044, -13811, -10566, -4400, -1009, 4193, 8907, 12614, 17000, 19658, 
    23051, 24919, 28084, 28502, 30345, 32515, 29574, 29599, 27748, 26069, 
    22316, 20747, 18976, 14256, 9492, 4883, 1873, -2832, -7985, -12905, 
    -16429, -18835, -23701, -25638, -26780, -30492, -30380, -31118, -31577, 
    -29902, -28679, -25185, -23376, -21900, -16300, -14012, -9710, -6023, 59, 
    5140, 7226, 10890, 16463, 18836, 22070, 25594, 28053, 30599, 29175, 
    29577, 30672, 29352, 28726, 26531, 23508, 20854, 18012, 13573, 8395, 
    5280, 689, -4011, -6488, -13603, -15044, -18818, -21679, -24293, -29057, 
    -30179, -29207, -31274, -31272, -28184, -28682, -26377, -24508, -20309, 
    -17890, -14255, -9982, -7087, -2342, 3465, 8233, 11584, 15013, 19084, 
    20972, 24506, 26689, 29163, 30976, 29922, 30559, 28674, 28394, 26326, 
    23275, 21612, 17556, 15546, 9811, 6834, 1479, -1446, -7894, -12253, 
    -15574, -20334, -22161, -25006, -26589, -30193, -29075, -30923, -30535, 
    -30048, -30495, -26116, -25570, -20071, -18355, -12751, -11576, -5933, 
    -1244, 3638, 7773, 10894, 14125, 19149, 21323, 23620, 27946, 28686, 
    29864, 29719, 30512, 28422, 27952, 26104, 25283, 21048, 17589, 14678, 
    9778, 6026, 1007, -1343, -8041, -10210, -16247, -18576, -21893, -24681, 
    -27225, -27747, -30356, -31450, -29871, -29792, -28689, -27023, -25594, 
    -20754, -17926, -13534, -9684, -5383, -1857, 2485, 5714, 11078, 14490, 
    19450, 21411, 23561, 26473, 28664, 30270, 29477, 30999, 30870, 28695, 
    26337, 24831, 20646, 19134, 15861, 11271, 6307, 3393, -1129, -6291, 
    -10480, -15734, -17571, -22379, -23249, -26151, -27572, -30185, -31317, 
    -29770, -30348, -28458, -27245, -25080, -22435, -18494, -15076, -10684, 
    -6957, -2566, 1040, 5781, 11185, 14151, 18903, 22379, 24510, 27615, 
    28630, 30236, 31562, 30772, 29696, 29402, 27280, 25945, 21668, 18265, 
    15368, 10659, 7118, 2924, -171, -6929, -8809, -14283, -19068, -21069, 
    -23945, -25972, -28365, -30636, -31711, -30880, -31171, -28057, -27528, 
    -25669, -22833, -19139, -14948, -11911, -7527, -1628, 2305, 5182, 10899, 
    13912, 17038, 20310, 24717, 26107, 28851, 31469, 29474, 31326, 30596, 
    29099, 26494, 24926, 22918, 19058, 16358, 10909, 7981, 3335, -1297, 
    -5466, -10466, -13410, -17705, -20506, -24371, -26211, -29146, -29913, 
    -30983, -30761, -30237, -30860, -27153, -24474, -22688, -19961, -16923, 
    -11053, -8098, -2470, 773, 5132, 9999, 12571, 17614, 19158, 24346, 25101, 
    28581, 29440, 31592, 31133, 30575, 29313, 27548, 24519, 21908, 20781, 
    14746, 10969, 8206, 5484, -1114, -4609, -8685, -14115, -16140, -20478, 
    -23583, -26853, -28337, -29554, -31275, -30871, -30406, -28779, -28101, 
    -26406, -23874, -20539, -17158, -12138, -9481, -3880, 592, 3395, 9297, 
    13301, 16172, 19901, 22980, 27499, 27709, 30241, 30050, 29136, 29817, 
    28075, 28789, 26206, 23319, 20171, 15665, 12164, 10003, 2330, -255, 
    -5439, -8262, -13649, -17303, -20381, -23842, -26589, -27199, -28520, 
    -31980, -30401, -30712, -28904, -28051, -25865, -24095, -20820, -16153, 
    -12604, -8459, -4300, 218, 3838, 9119, 14008, 16275, 18910, 24460, 26787, 
    27931, 29991, 29349, 29665, 31387, 28985, 29150, 25930, 23652, 20975, 
    16429, 12430, 9447, 4524, -521, -4894, -8854, -14431, -15218, -20099, 
    -23120, -25394, -27945, -29449, -29573, -30344, -29817, -30100, -29420, 
    -25869, -21786, -20572, -15642, -14136, -9969, -4684, -99, 4117, 9278, 
    12763, 16097, 21395, 21754, 24621, 27607, 28777, 29789, 29406, 28811, 
    30366, 27592, 26782, 24538, 19693, 18138, 13693, 10290, 5250, 1407, 
    -3477, -8159, -12058, -17401, -19453, -21721, -25685, -28441, -29822, 
    -31481, -30249, -29943, -29253, -29446, -26550, -23459, -21236, -17893, 
    -14578, -8696, -4027, -1040, 4248, 6584, 10774, 15905, 19369, 22197, 
    24565, 27790, 28534, 29862, 31075, 30062, 29445, 27925, 25970, 24190, 
    21936, 17379, 13194, 8107, 4843, 304, -3724, -7581, -11037, -15262, 
    -18122, -23522, -24204, -27095, -29179, -29664, -29358, -31575, -29952, 
    -28251, -27756, -24299, -20513, -17757, -13939, -10000, -7077, -1576, 
    3055, 7438, 12969, 15350, 17714, 21676, 25379, 28037, 30447, 32031, 
    31356, 30564, 29989, 27606, 26550, 23932, 21361, 16865, 13763, 10919, 
    7703, 1309, -1374, -8598, -9871, -15253, -17994, -22187, -25817, -28267, 
    -29046, -29071, -30187, -30582, -30236, -29613, -26295, -24249, -21043, 
    -18495, -13092, -8595, -7251, -2668, 3814, 6895, 10570, 14142, 17018, 
    21120, 23524, 27594, 29933, 30535, 31653, 30381, 29973, 29327, 27307, 
    24486, 22830, 18101, 16124, 10708, 5123, 3362, -2311, -5784, -9988, 
    -14121, -18239, -22821, -24711, -26753, -29455, -29964, -30912, -31394, 
    -30324, -28625, -27291, -25144, -22044, -16998, -14912, -10446, -6961, 
    -1722, 1951, 6104, 11768, 14195, 19229, 23041, 24891, 26069, 28618, 
    31759, 30893, 29570, 30159, 28838, 27676, 23756, 20374, 19403, 16542, 
    10832, 6222, 3522, -1094, -5558, -9574, -13552, -16682, -21373, -23033, 
    -27761, -29843, -28196, -31846, -31489, -29116, -28988, -26847, -24433, 
    -23153, -18665, -16198, -12416, -7344, -3085, 1401, 5950, 9758, 13508, 
    19232, 21778, 23015, 25582, 30275, 29398, 29475, 30798, 30540, 29473, 
    28321, 23820, 23268, 19245, 15650, 10186, 8137, 2771, -2753, -6543, 
    -11538, -13874, -17507, -19502, -22797, -26534, -28485, -31542, -30764, 
    -31649, -28991, -29692, -28245, -24956, -20926, -19704, -15596, -13481, 
    -8174, -1806, 1301, 6039, 10486, 13159, 17320, 20452, 25393, 26580, 
    28524, 29690, 30812, 29828, 30161, 28993, 27308, 25789, 23310, 19131, 
    15113, 12149, 6542, 3518, -371, -5693, -10534, -14118, -18055, -20490, 
    -24105, -25425, -30193, -29853, -30333, -29191, -29398, -29683, -27551, 
    -25737, -21408, -21033, -14260, -10904, -8287, -2879, -267, 5136, 9410, 
    14114, 17561, 20244, 24894, 27068, 27062, 29489, 30714, 30770, 30358, 
    29248, 27479, 24169, 21857, 20149, 15771, 13594, 7634, 4709, -1718, 
    -4894, -9671, -12556, -17507, -19809, -23857, -26146, -29242, -29853, 
    -30536, -31158, -30685, -29121, -28833, -24958, -22073, -19321, -16995, 
    -12401, -8401, -4044, 826, 5004, 8589, 13524, 15972, 20816, 25089, 25237, 
    28322, 28871, 31557, 29770, 31674, 29819, 27776, 26006, 23349, 20981, 
    15277, 12883, 8527, 4203, -29, -4456, -8511, -13530, -16309, -19508, 
    -22723, -24483, -27746, -28208, -31241, -31006, -30610, -29179, -28779, 
    -25352, -23411, -19936, -16381, -11917, -8631, -4318, 32, 4041, 9947, 
    14156, 17359, 20276, 24305, 25482, 29420, 29612, 30698, 31230, 30294, 
    28947, 27699, 26801, 24447, 19319, 16923, 13433, 8258, 4559, 316, -2906, 
    -7148, -13420, -18045, -19754, -22876, -26857, -27334, -29805, -29464, 
    -30549, -31070, -30390, -27073, -26468, -23511, -21175, -16275, -12497, 
    -10339, -3339, -26, 2110, 8061, 11973, 14751, 18537, 22497, 26468, 29279, 
    29329, 31718, 30523, 31479, 29801, 29314, 26725, 24077, 20559, 18539, 
    13255, 8600, 4735, 407, -3110, -6834, -12344, -16242, -20572, -22333, 
    -24615, -27119, -29559, -30719, -31232, -31711, -29538, -29471, -27143, 
    -24781, -20392, -16890, -12722, -10728, -5030, -1374, 4832, 7738, 12338, 
    14962, 18237, 21813, 26177, 27488, 28714, 29936, 31189, 29479, 28770, 
    27132, 26942, 23249, 22701, 18404, 13394, 8537, 4896, 1509, -3339, -7255, 
    -12759, -14701, -18250, -21435, -25172, -26055, -29727, -29732, -29819, 
    -29853, -28692, -30002, -26530, -23673, -22548, -17914, -13085, -9559, 
    -4295, -1617, 4146, 8048, 12746, 17075, 19349, 22781, 26475, 26562, 
    28575, 30447, 30565, 31663, 30486, 28589, 27366, 24426, 20176, 18720, 
    14243, 9947, 6853, 1270, -2406, -6198, -10738, -15279, -19718, -22047, 
    -25346, -27732, -30460, -30548, -32037, -30612, -31112, -28611, -27534, 
    -24206, -22039, -18163, -15054, -10536, -7232, -912, 1067, 5319, 12240, 
    15648, 19141, 21959, 25543, 25945, 28326, 30722, 30171, 29680, 31247, 
    29347, 27847, 24530, 20829, 18878, 15255, 9151, 6251, 3016, -1415, -7491, 
    -11102, -13917, -18548, -23345, -24014, -26189, -30593, -30164, -31731, 
    -32250, -29888, -29881, -27148, -24787, -21924, -17698, -14800, -11509, 
    -5173, -3600, 798, 7301, 10635, 15144, 19407, 22691, 23418, 27192, 29839, 
    29901, 30093, 30392, 31133, 28915, 26888, 23053, 21556, 19924, 14170, 
    11349, 5634, 1257, -2104, -6119, -9953, -14659, -18069, -20044, -23637, 
    -27237, -28896, -29878, -29372, -29505, -30091, -30562, -26697, -24912, 
    -20613, -18485, -14915, -10722, -5591, -871, 1510, 6034, 11154, 14699, 
    17695, 20132, 25097, 26999, 29136, 29849, 30631, 29952, 30062, 30232, 
    27699, 25768, 22363, 18785, 15471, 11473, 5658, 1688, -1795, -4901, 
    -8831, -14999, -18057, -20544, -24461, -25526, -27770, -29621, -29677, 
    -31000, -30589, -28968, -27022, -24630, -22366, -19697, -15213, -11591, 
    -7123, -2520, 2059, 6589, 8954, 13765, 17442, 20752, 23741, 27229, 28972, 
    29890, 31524, 30162, 31150, 29068, 28164, 24642, 22434, 17594, 15030, 
    11543, 7475, 3770, -479, -4455, -9877, -13095, -17451, -20855, -23106, 
    -24894, -27696, -28616, -31923, -30503, -29689, -29036, -26107, -24452, 
    -21054, -19341, -15698, -12425, -8114, -3093, -473, 4803, 10279, 13432, 
    18231, 20554, 24189, 25047, 27619, 28811, 30685, 29067, 29977, 28182, 
    27861, 25859, 21535, 20836, 17319, 12216, 8796, 4201, -622, -5312, -9586, 
    -13524, -15617, -19831, -25256, -26133, -28021, -28459, -32448, -31146, 
    -29317, -29315, -26891, -25759, -23284, -20253, -16125, -12175, -7879, 
    -2969, -151, 3370, 8364, 13323, 17191, 21657, 23229, 25853, 28530, 28362, 
    30240, 30517, 30572, 29618, 26791, 26800, 22884, 18431, 15192, 13607, 
    9200, 3796, 324, -4685, -8549, -14084, -16028, -19333, -23823, -26924, 
    -28202, -30846, -29524, -31259, -29944, -29934, -28082, -25878, -23424, 
    -21036, -17979, -12799, -8450, -4604, 774, 4163, 9381, 11916, 17693, 
    19269, 22435, 24658, 28157, 30394, 30402, 29897, 31768, 30420, 27529, 
    25610, 23887, 20783, 15841, 13650, 9100, 4171, 1366, -5369, -8115, 
    -12521, -16844, -19054, -22331, -26118, -27631, -28042, -28772, -30121, 
    -29923, -28398, -29057, -25291, -23814, -19143, -15306, -12381, -9032, 
    -5450, -412, 3930, 7369, 12222, 18152, 19241, 23022, 25843, 26589, 29663, 
    30643, 30483, 30551, 29507, 29090, 24421, 23847, 21448, 17665, 13770, 
    10203, 3928, 613, -3771, -7509, -11803, -15573, -19601, -21829, -26594, 
    -27848, -28780, -29594, -30320, -31108, -29470, -27493, -25608, -24360, 
    -20272, -17087, -12329, -8727, -4893, -1585, 3102, 7274, 13338, 15838, 
    20179, 22148, 25495, 27994, 27507, 30370, 32108, 30766, 30170, 28109, 
    26276, 23448, 19562, 17761, 14353, 9620, 6009, -662, -1738, -7285, 
    -12264, -16159, -20230, -21918, -26903, -27494, -28319, -31531, -30866, 
    -29432, -30287, -29115, -28044, -24285, -21043, -17667, -13434, -9726, 
    -3948, -691, 2489, 6677, 13205, 16091, 20301, 22350, 26302, 26965, 27544, 
    31081, 30983, 31896, 28496, 29249, 25723, 23734, 20394, 16979, 13582, 
    9058, 5152, 1701, -3323, -7424, -10068, -15179, -17071, -22249, -25100, 
    -27450, -27547, -29456, -30520, -31226, -31194, -28795, -26530, -24362, 
    -21318, -18166, -14322, -9349, -7374, -3069, 1403, 6200, 10881, 15730, 
    19977, 21048, 24756, 27430, 28943, 30223, 30716, 30952, 30449, 27880, 
    26153, 24600, 21834, 18655, 15549, 11854, 5937, 2319, -2312, -7871, 
    -11722, -15737, -19337, -22572, -24966, -26766, -29273, -30620, -29666, 
    -31160, -29618, -29070, -28543, -25737, -21437, -17293, -14295, -10050, 
    -4874, -2075, 3073, 7754, 10235, 15175, 17875, 22889, 25078, 26082, 
    28942, 30164, 29504, 29731, 29586, 27316, 25526, 24753, 21738, 19103, 
    14537, 11766, 7315, 2481, -1352, -5659, -10175, -12693, -19346, -21320, 
    -25255, -26825, -29153, -29439, -30715, -31481, -29941, -28034, -25866, 
    -25367, -23863, -18199, -14720, -10461, -5294, -2931, 2101, 6480, 9603, 
    14499, 18362, 22461, 25438, 28371, 28747, 31078, 30176, 31835, 30957, 
    30234, 28850, 25061, 22873, 18975, 15743, 10400, 8036, 2594, -2384, 
    -6136, -11971, -15296, -17494, -20520, -24958, -26289, -28498, -31341, 
    -31237, -30632, -30544, -29094, -28038, -25536, -21672, -18319, -16995, 
    -12501, -7138, -2356, 2498, 5519, 10347, 12909, 18923, 21481, 25084, 
    27072, 27288, 29209, 30304, 31470, 31733, 29671, 27114, 25603, 21823, 
    20555, 16647, 10869, 7682, 3820, -1486, -5510, -10430, -13957, -18512, 
    -19512, -23232, -26253, -28114, -28520, -31148, -29871, -30787, -29854, 
    -28277, -24428, -22537, -21074, -15204, -11451, -8464, -3685, 291, 5048, 
    9414, 13550, 18513, 20265, 23203, 25089, 30044, 28241, 29317, 30878, 
    30515, 28632, 28218, 26097, 22653, 18713, 17051, 12870, 9184, 5361, 286, 
    -4995, -9880, -13563, -16590, -20832, -23686, -26148, -28484, -28648, 
    -30728, -30632, -30685, -28959, -28172, -26616, -24595, -18912, -16435, 
    -13727, -7518, -3305, 584, 4399, 8880, 12294, 17620, 20335, 25065, 24707, 
    28231, 28814, 29329, 30095, 30329, 30094, 27170, 25861, 24854, 20548, 
    16966, 13141, 7238, 3201, -841, -5994, -7592, -12888, -17875, -19085, 
    -21679, -25992, -28458, -29654, -30998, -30447, -31075, -29535, -27901, 
    -26835, -23909, -19595, -16895, -12406, -9723, -2842, -819, 5674, 9466, 
    13224, 17863, 18806, 22428, 26093, 28025, 29193, 29599, 31767, 31415, 
    30399, 28271, 25228, 24384, 19828, 15963, 13178, 9259, 5858, 122, -3825, 
    -7322, -11670, -14904, -19445, -23200, -25197, -28356, -29983, -30747, 
    -31008, -30380, -29519, -28569, -25331, -24344, -20491, -17394, -13746, 
    -7916, -6309, -1309, 3251, 9398, 12581, 15267, 19742, 23971, 27260, 
    26824, 29362, 30274, 31858, 31300, 29665, 27935, 26463, 23945, 21481, 
    15911, 12873, 9240, 4935, 757, -3316, -8051, -12366, -15912, -19732, 
    -23403, -25796, -27689, -29590, -29851, -31163, -31587, -29972, -27293, 
    -26199, -24626, -22222, -17910, -13649, -9722, -6035, 831, 3889, 8621, 
    11329, 14418, 19784, 23074, 25461, 25975, 28798, 29775, 31284, 30214, 
    30018, 28131, 26439, 25289, 20899, 17428, 13394, 9677, 5441, 1725, -3794, 
    -6829, -10725, -16340, -20171, -22565, -24452, -27280, -29525, -29193, 
    -30128, -32195, -30261, -28282, -26510, -25301, -21419, -16554, -13529, 
    -11007, -4109, -1748, 3626, 6679, 11713, 14948, 18553, 23384, 25905, 
    27432, 29565, 29502, 29539, 30207, 31437, 27960, 26300, 24922, 21634, 
    17750, 13728, 9990, 7041, 1274, -3979, -7921, -12096, -15520, -18087, 
    -23106, -24420, -26023, -30020, -29146, -31167, -32169, -29554, -29172, 
    -25334, -24533, -21471, -18714, -15229, -10610, -5136, -3052, 3017, 7897, 
    11400, 15006, 18845, 21178, 24699, 28003, 29238, 30258, 29512, 29862, 
    30973, 30280, 27055, 24862, 21499, 17863, 14526, 9997, 6203, 901, -1557, 
    -5254, -11330, -14401, -18656, -21244, -24657, -27858, -29085, -30448, 
    -32170, -30706, -30770, -29195, -27435, -24105, -22346, -17553, -14516, 
    -10032, -5578, -2602, 2485, 6638, 10692, 14246, 18562, 22181, 24351, 
    26724, 28871, 30142, 32100, 30222, 29254, 28433, 26598, 25438, 21509, 
    19421, 13684, 10968, 5616, 2749, -2929, -6137, -10051, -13796, -18896, 
    -22466, -24968, -25903, -29344, -29762, -30308, -31252, -29436, -28147, 
    -28010, -24237, -22594, -19685, -14495, -9712, -6940, -1486, 1061, 7054, 
    11536, 14398, 17728, 21003, 23521, 25900, 28825, 29724, 30326, 30478, 
    28755, 27445, 27944, 25355, 22683, 19230, 15045, 12290, 7595, 2650, 
    -2373, -4956, -11145, -13068, -17451, -20561, -23866, -25932, -27897, 
    -29326, -31082, -29528, -30254, -27761, -27061, -24728, -21825, -20794, 
    -16170, -11624, -8025, -2751, 2399, 5432, 10175, 13499, 17208, 20894, 
    23773, 25837, 27981, 28969, 30193, 30965, 31556, 27834, 27509, 25175, 
    24295, 20743, 15234, 11553, 6982, 4033, -551, -3985, -9779, -13224, 
    -17045, -19900, -22749, -25673, -28002, -31516, -30607, -29243, -31116, 
    -27743, -28731, -24634, -23656, -20635, -15339, -12651, -9359, -4540, 
    903, 7031, 8765, 13273, 18930, 21912, 24202, 26854, 28326, 29486, 30214, 
    29837, 30791, 28351, 26239, 26426, 23586, 19807, 15276, 11906, 6900, 
    4166, -179, -3595, -10243, -12711, -17747, -21264, -22785, -25638, 
    -27970, -30041, -31479, -31091, -30923, -30072, -27480, -26320, -21677, 
    -21002, -17453, -12019, -8375, -3414, 372, 5504, 9020, 12397, 17790, 
    20267, 23313, 25008, 27367, 28549, 31604, 30917, 30773, 30190, 28600, 
    26323, 24705, 19066, 16164, 11452, 8740, 3209, -246, -4609, -8237, 
    -11466, -16511, -19829, -24227, -26881, -27988, -28800, -29922, -31934, 
    -30118, -30180, -27822, -26403, -22816, -20319, -17984, -13429, -8694, 
    -3985, -855, 4598, 7302, 12885, 18405, 18855, 22378, 24771, 29505, 28143, 
    30423, 31627, 31643, 29046, 27467, 25631, 23849, 20512, 17863, 13514, 
    9442, 5027, -430, -5309, -8670, -13507, -16948, -19170, -22332, -25322, 
    -27761, -30163, -30669, -30331, -29748, -28044, -27602, -26607, -22600, 
    -20355, -16330, -12096, -8506, -3792, -1945, 4391, 8663, 12415, 14392, 
    19789, 22490, 26020, 27768, 29951, 30673, 31808, 31021, 30017, 29343, 
    26299, 23059, 21421, 17793, 13123, 9969, 3907, -170, -2815, -8922, 
    -12535, -16258, -18567, -23204, -26009, -28482, -29527, -29257, -30580, 
    -31047, -30061, -27032, -25656, -23676, -21782, -18506, -13374, -10824, 
    -5838, -1778, 4508, 7375, 11657, 15783, 20355, 23045, 24087, 27824, 
    29842, 31611, 32335, 31006, 30896, 28559, 26689, 24106, 21491, 16615, 
    14088, 9641, 5756, 1770, -2729, -7905, -11044, -15953, -20207, -23170, 
    -26766, -27536, -29846, -29820, -29764, -31572, -30026, -28499, -27243, 
    -23696, -20214, -17056, -14962, -10887, -6392, -1682, 3001, 7765, 11468, 
    15699, 20123, 21701, 24912, 28736, 29355, 30137, 31312, 31091, 30293, 
    27649, 26007, 23830, 21683, 17707, 14499, 9771, 6081, 1428, -4002, -7780, 
    -10773, -15601, -17449, -21724, -25648, -27301, -29378, -30312, -30561, 
    -29628, -29447, -29069, -27045, -25085, -22160, -18050, -14823, -9334, 
    -6556, -2799, 2485, 7660, 11491, 14838, 19827, 21628, 24705, 28498, 
    29223, 30458, 29494, 30294, 29388, 28050, 26349, 24536, 22611, 18360, 
    15063, 10918, 6339, 773, -3712, -6493, -11406, -14795, -18562, -23261, 
    -24990, -26922, -29409, -29595, -31201, -31128, -31170, -27095, -25548, 
    -25859, -22591, -18044, -13802, -12247, -6848, -2003, 2199, 6593, 10231, 
    16328, 17770, 20761, 24117, 27164, 28235, 29962, 29381, 30770, 29346, 
    30080, 26430, 24475, 22430, 19950, 15291, 11649, 6483, 2794, -2328, 
    -6315, -11723, -13709, -18455, -21810, -24295, -28197, -28808, -29185, 
    -29524, -31642, -29576, -29320, -27722, -24523, -21892, -20418, -14808, 
    -10300, -6159, -1910, 1254, 5760, 8544, 14267, 17457, 21965, 24428, 
    27519, 27442, 29855, 29961, 31190, 30178, 28502, 26548, 25333, 23947, 
    20104, 16982, 12599, 6734, 2241, -1697, -7330, -11226, -14088, -17570, 
    -21268, -25255, -26380, -26895, -29657, -31401, -30059, -30431, -29281, 
    -25683, -23526, -23821, -19129, -14720, -10878, -7016, -3870, 1357, 5551, 
    10673, 14808, 17204, 21324, 23242, 27508, 28041, 29776, 30666, 31328, 
    29110, 29008, 27180, 23680, 21832, 19963, 15541, 12319, 6933, 3048, 374, 
    -5287, -10289, -13003, -17895, -19144, -23652, -26756, -28681, -29476, 
    -30496, -31061, -30395, -28986, -26581, -25409, -22323, -19909, -16224, 
    -10423, -7739, -3399, 1323, 4523, 9264, 14007, 16790, 19281, 23326, 
    27718, 26838, 29686, 30959, 32239, 30141, 29221, 27127, 25259, 24316, 
    21191, 16102, 12316, 7341, 4218, -485, -5506, -8888, -14541, -17566, 
    -19974, -23143, -24761, -27318, -28195, -31282, -32531, -30078, -29982, 
    -28443, -25567, -23804, -21102, -14858, -11970, -8677, -3600, 780, 5678, 
    10714, 14062, 17763, 21550, 23433, 26715, 28718, 29349, 31392, 32107, 
    31720, 30310, 28922, 25746, 23855, 18674, 16102, 11923, 8967, 4613, 
    -1052, -6156, -9665, -12853, -17580, -20067, -22294, -25469, -27826, 
    -30151, -29745, -30945, -30063, -28760, -29602, -26877, -23245, -20280, 
    -17635, -14028, -9209, -5706, 1467, 4754, 9487, 11832, 15504, 20131, 
    22283, 25622, 27521, 29246, 30273, 31280, 31452, 28686, 28241, 26013, 
    23715, 21831, 18481, 12359, 7554, 3421, -156, -3392, -7910, -12597, 
    -15404, -19939, -23503, -26614, -28553, -29202, -31560, -31143, -31329, 
    -30186, -26889, -25645, -23567, -21328, -17478, -13526, -9146, -4054, 
    255, 5244, 8605, 12175, 16073, 20468, 23973, 26364, 27259, 29080, 31519, 
    31023, 30289, 30534, 28037, 25519, 23195, 21050, 17177, 12574, 8496, 
    3979, 941, -4775, -9199, -12961, -14620, -19735, -22963, -25464, -28393, 
    -28936, -29887, -31299, -30300, -30280, -27978, -25257, -22430, -20646, 
    -16677, -13154, -8636, -4814, -806, 3765, 6596, 11608, 17559, 19545, 
    21537, 23613, 25917, 29673, 30638, 29819, 30426, 28921, 28924, 26891, 
    23801, 21656, 19078, 14297, 10128, 5473, 1495, -2348, -8690, -11592, 
    -15620, -19040, -22481, -26130, -26700, -28388, -30323, -29780, -29967, 
    -28666, -29180, -25052, -22845, -21036, -17859, -13641, -8583, -6367, 
    -486, 2174, 7295, 12603, 14310, 20409, 22774, 23446, 27911, 30488, 29386, 
    30867, 30764, 29040, 28756, 26379, 25188, 21022, 16873, 14946, 9898, 
    5806, -76, -2561, -7791, -10951, -16496, -19104, -22369, -26027, -27591, 
    -29611, -29691, -30525, -32016, -29819, -28739, -27171, -22905, -22771, 
    -19274, -14274, -9594, -5424, -976, 3622, 7771, 12126, 14238, 17073, 
    21169, 24587, 28866, 30554, 30493, 29631, 31594, 30157, 27560, 27205, 
    24497, 22138, 19748, 15599, 10006, 5927, 1644, -2265, -6078, -11565, 
    -14419, -17795, -20630, -26107, -27239, -28247, -30304, -31441, -29475, 
    -29275, -28939, -26394, -23472, -22894, -18367, -15862, -9481, -5576, 
    -3190, 2310, 5201, 11052, 14855, 17781, 22693, 24446, 27104, 28913, 
    29973, 32027, 31040, 30442, 28109, 27101, 24945, 21411, 17506, 14876, 
    10951, 5899, 3126, -2123, -7290, -11582, -15293, -18621, -20418, -26056, 
    -26917, -29852, -29427, -30760, -30932, -29459, -28985, -27684, -24703, 
    -20866, -19730, -16421, -10953, -6881, -2572, 1916, 7156, 11467, 13793, 
    17272, 21583, 24654, 26889, 28456, 30311, 29350, 30706, 31296, 28209, 
    26782, 26415, 21252, 18050, 15939, 12302, 6314, 2649, -1063, -4435, 
    -10708, -14718, -18887, -20486, -23851, -27078, -27841, -28690, -30001, 
    -30819, -28800, -28085, -27275, -25009, -20791, -18244, -15085, -10369, 
    -7627, -2848, 470, 6408, 11505, 13008, 19087, 20344, 24460, 27552, 29563, 
    29851, 31025, 31156, 29531, 30014, 26249, 25302, 20806, 20262, 15515, 
    13043, 7260, 4755, -945, -6188, -10730, -12489, -17741, -21669, -25521, 
    -25841, -28538, -28419, -31578, -30708, -30770, -29016, -27301, -26312, 
    -22481, -19677, -16546, -12236, -6554, -3090, 1979, 5786, 9441, 12780, 
    16576, 20108, 23353, 25777, 29087, 31130, 30796, 30761, 30431, 29417, 
    26443, 25512, 23676, 19405, 15750, 11390, 8790, 4774, -42, -5486, -8769, 
    -12055, -16963, -22192, -24301, -25700, -30105, -28292, -31090, -31961, 
    -32017, -30518, -27581, -24266, -22699, -18959, -14566, -11151, -9460, 
    -4684, 353, 3672, 9226, 14959, 16166, 20210, 23215, 27072, 28559, 31248, 
    30725, 29907, 31205, 30209, 26532, 25661, 23781, 19853, 16150, 11930, 
    8904, 3960, -617, -4956, -8494, -12642, -16383, -21242, -23031, -25206, 
    -27190, -28470, -29490, -30784, -30441, -29898, -27603, -26142, -22754, 
    -19811, -16800, -13115, -9085, -3226, -245, 4287, 8061, 12091, 15455, 
    19261, 24133, 25693, 26386, 29214, 31680, 30832, 31130, 30551, 28484, 
    27179, 23785, 20082, 16692, 12798, 8864, 4715, 488, -3957, -8512, -11618, 
    -17578, -19129, -23989, -24702, -27742, -31234, -30235, -31273, -31781, 
    -28035, -29001, -24527, -22948, -19830, -15711, -12614, -10175, -4251, 
    -504, 4162, 8732, 11073, 15810, 19566, 23626, 26834, 28961, 28951, 31095, 
    31142, 31518, 28404, 29477, 26354, 23867, 20543, 16569, 13784, 10230, 
    5315, 1412, -3616, -8720, -11225, -16384, -19887, -23121, -24805, -27549, 
    -29474, -31063, -29792, -29514, -29086, -28803, -25912, -25301, -19413, 
    -16275, -14889, -8398, -4440, -175, 3377, 6208, 11602, 16954, 19457, 
    23170, 25551, 28289, 30140, 29975, 30445, 29340, 30334, 27455, 27301, 
    23628, 21295, 16324, 14225, 9468, 5818, 1717, -2616, -7451, -12181, 
    -15329, -18804, -22220, -25347, -28011, -28741, -29866, -30929, -29910, 
    -28982, -28703, -27293, -23143, -21428, -17600, -14008, -8604, -4424, 
    -547, 2741, 6788, 11352, 16945, 18682, 22553, 26040, 27668, 28284, 31639, 
    30663, 31771, 30710, 30065, 25252, 23493, 21104, 19510, 14288, 9571, 
    5707, 694, -1256, -8793, -9714, -15185, -19603, -22174, -24825, -27205, 
    -28931, -31060, -30897, -30949, -29673, -27335, -26296, -24245, -21683, 
    -18288, -14155, -10543, -6528, -1582, 2392, 5946, 10671, 13570, 19487, 
    21531, 25436, 26115, 29854, 30244, 31994, 31352, 31208, 28128, 26337, 
    25645, 21909, 18304, 15775, 9798, 6889, 2890, -2095, -7092, -11471, 
    -14757, -17105, -22528, -24202, -26971, -29814, -29107, -30585, -30869, 
    -28629, -30519, -27908, -23891, -21211, -18440, -14500, -10605, -7148, 
    -1466, 3828, 6503, 10945, 14995, 19372, 22951, 24333, 27543, 28080, 
    29943, 30301, 31221, 30687, 28891, 27956, 24744, 21108, 17523, 14672, 
    10502, 6475, 3720, -3323, -4976, -9254, -15068, -17327, -21522, -25377, 
    -26887, -29242, -31393, -29645, -31369, -30163, -28959, -26423, -25098, 
    -21602, -18243, -13981, -9888, -7138, -2501, 1725, 7170, 10557, 13003, 
    18964, 21760, 23215, 28086, 28758, 30505, 31528, 30967, 30117, 30449, 
    27863, 25374, 22819, 19260, 16534, 11615, 8524, 3770, -2326, -4659, 
    -9560, -14300, -17240, -20524, -24308, -26493, -27700, -29126, -30793, 
    -31578, -30061, -28898, -28678, -24320, -22734, -18968, -14629, -13023, 
    -7110, -3842, 517, 4199, 10059, 14033, 17704, 22698, 24233, 26256, 28968, 
    29937, 30641, 31455, 31208, 28763, 26910, 25963, 21430, 18728, 14438, 
    12613, 8075, 3156, 253, -5544, -10174, -14884, -18049, -21143, -24054, 
    -26080, -29439, -28963, -30979, -32232, -31774, -30785, -27273, -24852, 
    -22935, -20623, -15658, -11952, -7118, -4472, -574, 4215, 11030, 13386, 
    16850, 20588, 22785, 26779, 30252, 30508, 30886, 29420, 30648, 30001, 
    29355, 25541, 21603, 19009, 15070, 11971, 7755, 3178, -2070, -4283, 
    -8373, -13589, -15656, -20913, -23037, -25991, -28560, -30704, -30555, 
    -30624, -30076, -29809, -26720, -25473, -23530, -20015, -15822, -12925, 
    -8762, -4707, 306, 5458, 8625, 13655, 18086, 20913, 23853, 26475, 28012, 
    30704, 29549, 31046, 29406, 31292, 27157, 26119, 22789, 20097, 15712, 
    13939, 8616, 3600, -1392, -3073, -9568, -13469, -16843, -21111, -23229, 
    -26437, -26656, -30735, -31248, -31573, -30173, -30517, -27331, -25088, 
    -22197, -19086, -16255, -13482, -8079, -4277, -541, 3823, 8900, 13481, 
    15832, 21092, 22906, 26823, 27616, 30262, 30409, 30035, 29910, 30168, 
    26535, 24884, 24665, 21028, 17681, 11468, 8262, 5287, -370, -2906, -7334, 
    -12967, -17101, -19507, -23266, -25832, -27656, -29860, -30740, -31679, 
    -30378, -30821, -29032, -25948, -24319, -20082, -17967, -12939, -10272, 
    -4832, -1601, 4224, 8719, 13365, 16269, 20378, 23206, 24702, 28919, 
    28927, 30451, 31876, 30754, 29610, 29329, 25306, 24281, 21539, 17909, 
    13390, 8229, 6508, -703, -3119, -8571, -11083, -15857, -21113, -21785, 
    -25459, -27291, -29926, -31343, -31287, -30541, -27887, -27894, -25666, 
    -23713, -21235, -17871, -13639, -9970, -5106, -1421, 4264, 8229, 11224, 
    15048, 19571, 23515, 25939, 27816, 30530, 31371, 30937, 30682, 29017, 
    27489, 26422, 22458, 19347, 17513, 12785, 9183, 4591, 61, -3392, -6741, 
    -12992, -16637, -18291, -23168, -24898, -26373, -29030, -29705, -29407, 
    -29301, -28379, -28680, -27235, -24653, -20688, -16978, -14944, -8875, 
    -6312, -2402, 2717, 7281, 13051, 15369, 18308, 22762, 25348, 28925, 
    29089, 29196, 29886, 32060, 30234, 28186, 27153, 25815, 22497, 18232, 
    15117, 9562, 6809, 1592, -2339, -6053, -10893, -14123, -18020, -22412, 
    -23778, -27089, -28839, -30362, -30823, -31537, -30030, -28737, -26182, 
    -23588, -20920, -19351, -13500, -8647, -6367, -1515, 1640, 5272, 10033, 
    14434, 19628, 20382, 25152, 26733, 27481, 30639, 29417, 30245, 29493, 
    27871, 26266, 24959, 22349, 18364, 13408, 11453, 7745, 1075, -2396, 
    -7309, -12011, -14714, -17159, -23511, -23999, -27820, -28807, -30577, 
    -32287, -31051, -30935, -27636, -27394, -24358, -21987, -17922, -15693, 
    -10103, -8178, -895, 2216, 6314, 11531, 16648, 18504, 21971, 25692, 
    27039, 28400, 30099, 31131, 31672, 30232, 28655, 27668, 24715, 22441, 
    19904, 13458, 10491, 6979, 2772, -1626, -5893, -10686, -14843, -19006, 
    -21401, -24680, -26215, -28657, -29026, -30576, -30646, -29590, -29535, 
    -27421, -24766, -21081, -17764, -15576, -10942, -7074, -1467, 2033, 6441, 
    9586, 15232, 19060, 21141, 23450, 27123, 28726, 28927, 32148, 30574, 
    30186, 28885, 27724, 25223, 22165, 19616, 15824, 12435, 6852, 3760, 
    -1525, -5774, -11511, -12791, -19267, -21329, -25369, -26652, -29393, 
    -31057, -31047, -31614, -29309, -28516, -28359, -24999, -22293, -18979, 
    -16051, -11753, -7852, -2849, 1591, 5590, 8982, 14158, 18229, 21705, 
    24117, 26496, 28955, 30885, 30879, 31916, 29360, 28824, 27368, 25918, 
    23288, 19076, 14800, 12368, 5870, 2510, -1729, -4854, -8231, -15179, 
    -17740, -21761, -23894, -26806, -27025, -29182, -29458, -29517, -31466, 
    -29403, -26984, -24885, -21599, -19567, -15555, -10841, -9266, -3781, 
    620, 5484, 10198, 12689, 18121, 20511, 24090, 27466, 28538, 29342, 30396, 
    31054, 31665, 29992, 26222, 25124, 24310, 20617, 16350, 12251, 9101, 
    3095, -1030, -4132, -9797, -12844, -16932, -19166, -24430, -26061, 
    -28175, -28761, -31210, -31864, -31173, -30205, -27657, -25512, -23420, 
    -20671, -16612, -11179, -8452, -3014, -267, 3152, 9369, 12730, 18417, 
    20861, 24506, 25505, 26557, 30932, 29634, 29850, 30561, 30145, 27892, 
    26914, 22123, 18901, 16684, 12750, 6985, 3356, 1121, -3733, -8567, 
    -11608, -15276, -21068, -24661, -24723, -29214, -29442, -30252, -29595, 
    -30931, -30288, -26588, -25509, -22696, -20687, -15419, -14275, -9724, 
    -4568, -353, 5338, 7462, 12107, 18053, 20221, 23432, 26317, 27769, 30094, 
    29664, 30916, 29163, 29411, 29242, 26144, 22901, 21161, 17275, 14271, 
    8098, 3977, -1261, -3328, -9280, -13013, -16423, -20693, -22886, -25632, 
    -27011, -28514, -31234, -31267, -31431, -29330, -29605, -27536, -22419, 
    -19552, -17219, -12563, -8576, -4073, -2012, 3559, 7325, 12903, 16373, 
    18779, 23103, 25519, 26749, 29823, 31700, 31369, 30728, 28198, 28595, 
    26003, 23342, 20310, 16064, 13646, 9220, 5395, 2093, -3014, -7954, 
    -13028, -15679, -18765, -21692, -24616, -28203, -28574, -29396, -29692, 
    -30648, -28704, -29618, -25807, -22506, -21585, -17128, -13369, -9223, 
    -4707, -806, 3078, 8291, 11815, 15756, 19778, 23079, 24743, 26568, 28864, 
    30739, 29714, 30579, 30412, 27642, 25959, 24472, 20037, 17628, 13920, 
    9620, 6174, 1711, -2764, -8218, -12919, -16085, -18568, -22424, -24746, 
    -27861, -28249, -29793, -31263, -31156, -29464, -29257, -25220, -24700, 
    -21323, -16478, -12851, -11532, -4496, -1311, 2832, 6134, 11406, 15988, 
    19619, 22619, 23944, 27805, 27846, 30098, 30293, 30902, 30675, 28969, 
    26674, 23586, 20552, 19519, 14233, 9315, 4786, 1851, -2352, -7012, 
    -11133, -13886, -17608, -22067, -25821, -27517, -28903, -30107, -31331, 
    -30465, -28858, -28999, -27907, -24363, -20940, -18243, -13160, -10090, 
    -7422, -2344, 2051, 6142, 9499, 15918, 18886, 22591, 24870, 26807, 29133, 
    30180, 29756, 31682, 30166, 29194, 26699, 23187, 21333, 19507, 14737, 
    10719, 6730, 1027, -3703, -6063, -11261, -13637, -19208, -22281, -24038, 
    -26461, -30197, -29185, -30902, -31272, -30948, -27479, -26117, -24115, 
    -20920, -17106, -14845, -11259, -7777, -2115, 2535, 6551, 9437, 14618, 
    17302, 22989, 24343, 27054, 28390, 28443, 32196, 30933, 30649, 29144, 
    26421, 23897, 21450, 18461, 13287, 10106, 7850, 1191, -2064, -6332, 
    -11012, -14650, -17358, -21428, -23829, -27136, -30004, -30243, -30480, 
    -30814, -30501, -28075, -28627, -24654, -22924, -19217, -15560, -11841, 
    -8085, -1919, 2650, 6758, 10463, 14022, 17949, 21919, 24533, 26734, 
    27051, 30520, 30766, 30211, 31866, 29903, 27665, 24652, 21332, 18829, 
    15231, 11877, 6305, 2837, -1005, -6857, -9198, -15402, -17053, -20695, 
    -24907, -27399, -28723, -29011, -30244, -30141, -30399, -30460, -27367, 
    -23839, -21440, -19607, -17021, -11265, -8328, -2527, 561, 5339, 9239, 
    15228, 17369, 21866, 25261, 27192, 28747, 29769, 31559, 29971, 28452, 
    28415, 26956, 24364, 22122, 18783, 15499, 13233, 8241, 3490, -673, -5999, 
    -9288, -14562, -16230, -20977, -23401, -24952, -28208, -29570, -30685, 
    -30280, -30386, -28463, -28705, -24000, -23138, -20971, -14991, -10678, 
    -7327, -3028, 865, 5341, 10619, 14321, 16595, 21883, 25539, 25354, 29424, 
    31036, 30363, 30239, 31636, 28109, 27754, 25023, 22592, 19435, 15216, 
    13587, 7702, 3489, -141, -5146, -7931, -14430, -17376, -22196, -23207, 
    -26125, -29286, -29579, -29874, -30825, -29924, -29787, -26874, -26177, 
    -22024, -19845, -16918, -12486, -8501, -4026, 1314, 5490, 8770, 13273, 
    16100, 18991, 24602, 25105, 28351, 29232, 29744, 30823, 30202, 29631, 
    26914, 26557, 21403, 19960, 16412, 11860, 8809, 5466, -262, -3160, -9189, 
    -11278, -16250, -21165, -22534, -26002, -27779, -29299, -30904, -30949, 
    -29553, -29579, -28443, -26756, -23649, -20514, -17335, -12631, -8611, 
    -5500, 418, 4522, 8634, 12830, 16124, 18835, 22489, 26791, 28925, 28236, 
    30379, 31009, 30653, 30796, 27891, 27031, 22775, 19962, 16288, 12978, 
    8589, 5539, 789, -4933, -8211, -13356, -16395, -19639, -22353, -24018, 
    -28519, -29472, -30412, -30908, -30829, -29175, -26718, -26252, -25122, 
    -20223, -18430, -12797, -10321, -5154, -1274, 5028, 8016, 12736, 16526, 
    20565, 23990, 25963, 29269, 30151, 29662, 30742, 30804, 29948, 30117, 
    26240, 24162, 19432, 16506, 14476, 10415, 5433, -171, -5144, -6441, 
    -10822, -16920, -21211, -23630, -24490, -28767, -29644, -28929, -30147, 
    -30902, -30081, -29139, -26936, -24743, -22118, -18062, -13623, -9970, 
    -5013, -357, 5137, 8359, 11418, 16095, 20688, 22701, 27178, 25963, 27995, 
    29569, 29356, 29818, 30763, 29567, 26883, 24846, 22108, 16482, 12044, 
    9746, 4647, 1837, -3627, -7913, -12233, -14361, -18966, -23132, -25962, 
    -27345, -30899, -32034, -29770, -31178, -30369, -28766, -27047, -24360, 
    -21422, -17711, -14300, -11111, -6860, 33, 3342, 7527, 11061, 17276, 
    18357, 23436, 26214, 26979, 28948, 30411, 31612, 31930, 29098, 28562, 
    27460, 24297, 20849, 17813, 14292, 10488, 5750, 1582, -3702, -8231, 
    -11537, -14753, -18604, -23305, -24672, -26525, -29337, -30596, -29673, 
    -30936, -31279, -28740, -25209, -24437, -21291, -17295, -14530, -11300, 
    -6207, -2186, 873, 5714, 12459, 14807, 18249, 21427, 24853, 27232, 28571, 
    31879, 31851, 30237, 28480, 27563, 26382, 23963, 21398, 18532, 14278, 
    11685, 5601, 1671, -1297, -7379, -10001, -15094, -19298, -23212, -24300, 
    -26593, -27540, -30094, -30047, -31134, -30715, -30311, -25336, -23484, 
    -21913, -18248, -15072, -10784, -6184, -2853, 3606, 6972, 9366, 14995, 
    17396, 19877, 25728, 28328, 27282, 29722, 30722, 30837, 29870, 30129, 
    25537, 24664, 20962, 18543, 14981, 11273, 5504, 2910, -1748, -7447, 
    -11378, -14440, -18344, -21615, -24840, -26765, -29028, -29886, -29478, 
    -30932, -28873, -29112, -26476, -25760, -21773, -17382, -14871, -11925, 
    -6655, -2433, 2086, 6659, 11550, 13687, 18748, 21782, 24744, 26745, 
    26901, 29428, 30031, 29819, 30638, 29853, 27604, 23509, 21276, 18700, 
    13463, 11227, 7268, 1954, -2116, -5043, -9829, -13824, -18272, -20539, 
    -25567, -26539, -29329, -30185, -29373, -30536, -30465, -29416, -26736, 
    -26147, -23295, -18702, -14500, -11357, -7425, -3736, -331, 5609, 9023, 
    14554, 17031, 21263, 24398, 26772, 28667, 30267, 30984, 30583, 28887, 
    27952, 26994, 25885, 21767, 19442, 15632, 12551, 6850, 4008, -1192, 
    -5525, -9375, -12798, -16908, -21562, -24592, -25646, -28868, -29795, 
    -29130, -30628, -29957, -29728, -27713, -24625, -21457, -18525, -14263, 
    -12059, -8040, -2386, 1296, 4369, 9658, 13876, 17170, 19672, 23291, 
    25774, 28812, 30216, 30029, 29592, 29252, 28951, 27552, 25849, 21931, 
    18914, 15559, 13655, 6949, 3958, -274, -4724, -8911, -14198, -17397, 
    -20626, -22796, -24444, -28926, -30167, -31552, -32296, -30319, -28303, 
    -27729, -25728, -22056, -20206, -16682, -12580, -8069, -4954, -149, 4734, 
    8278, 13978, 17236, 19839, 22629, 26173, 27279, 30428, 29731, 30775, 
    30686, 30079, 28655, 24908, 23226, 18405, 15107, 12124, 9658, 3934, 1414, 
    -4172, -9027, -11928, -17306, -18903, -22415, -26770, -28005, -30209, 
    -29264, -29669, -31158, -29133, -29163, -24862, -23550, -20229, -17771, 
    -12315, -7891, -4830, -1057, 3025, 9712, 12840, 18116, 19832, 24492, 
    27495, 28134, 29449, 29742, 30304, 29354, 29598, 28342, 26996, 22721, 
    21432, 15862, 13778, 8656, 5136, 1071, -3482, -7700, -12256, -15722, 
    -20525, -22231, -25759, -28450, -29392, -30529, -30251, -30961, -28998, 
    -28784, -26204, -22668, -20034, -16347, -13379, -8000, -5241, 231, 4258, 
    8557, 12712, 17158, 19837, 23760, 25734, 27886, 28665, 30883, 31966, 
    30717, 28839, 29802, 27137, 23732, 20712, 16422, 12116, 10052, 4990, 
    1772, -2956, -8099, -10913, -16937, -19153, -22961, -25158, -27995, 
    -29348, -31102, -31032, -29806, -30275, -29942, -26099, -24439, -20832, 
    -17924, -13227, -10758, -5789, -19, 4715, 7377, 10677, 16859, 18826, 
    22895, 25810, 26606, 29455, 29032, 30968, 31997, 29822, 29931, 26819, 
    24604, 21549, 18911, 13887, 9983, 3531, 8, -2776, -7471, -13421, -15191, 
    -19998, -23415, -24181, -29266, -28227, -31280, -32012, -30624, -30889, 
    -29982, -26123, -25456, -20856, -17788, -13339, -9022, -5073, -1269, 
    3212, 7170, 10167, 15604, 20470, 20952, 24388, 26905, 29853, 31831, 
    30290, 31374, 30499, 28757, 25561, 24502, 20056, 17515, 13659, 10616, 
    7378, 1931, -2688, -7860, -11196, -16824, -19595, -21028, -24242, -28426, 
    -29111, -30130, -30796, -31227, -30317, -29515, -27153, -24864, -20888, 
    -19490, -12814, -12181, -5692, -3125, 2130, 7087, 12539, 15377, 19124, 
    21568, 25272, 26605, 28525, 30217, 31280, 30841, 29187, 28658, 27566, 
    24805, 21688, 17620, 14545, 10368, 5997, 2170, -2167, -5958, -10645, 
    -14326, -19084, -22592, -24502, -27606, -29501, -29891, -29305, -30431, 
    -28298, -28588, -25901, -26102, -22458, -18849, -16083, -10492, -6173, 
    -512, 2160, 5594, 10088, 13468, 18362, 22935, 25147, 26472, 28244, 29729, 
    31559, 30828, 30476, 29223, 26478, 24225, 20424, 19506, 15404, 11167, 
    7733, 1034, -3013, -6759, -10237, -15296, -18534, -20498, -25679, -26442, 
    -28765, -31171, -31279, -30765, -29857, -29147, -25535, -25534, -20747, 
    -17624, -15814, -11805, -6950, -2698, 434, 5042, 11650, 15057, 17941, 
    20931, 24089, 27732, 27214, 30773, 30179, 30141, 29284, 29386, 26601, 
    25058, 22169, 19009, 15054, 11584, 7334, 3737, -769, -4640, -9189, 
    -13570, -17621, -21931, -24631, -25765, -28311, -28616, -30541, -30026, 
    -31382, -28285, -27323, -24883, -23202, -18193, -15196, -10766, -7146, 
    -2204, 1760, 4099, 11323, 14220, 17754, 21455, 23952, 27177, 27413, 
    29790, 30383, 31277, 29375, 29087, 26688, 25377, 22964, 19404, 15973, 
    11177, 7395, 3597, 39, -5775, -8825, -13327, -18681, -20250, -23021, 
    -25957, -28344, -28450, -30827, -30786, -30505, -29465, -26692, -26658, 
    -23960, -18758, -15706, -10959, -7643, -2579, 261, 5231, 9205, 13309, 
    17431, 21190, 24309, 25365, 26892, 29663, 30202, 31618, 30335, 28493, 
    28532, 24326, 21698, 19434, 15897, 12383, 8251, 3597, -644, -4358, -8642, 
    -12852, -18642, -21270, -24818, -25765, -27077, -29570, -31166, -30972, 
    -30650, -28960, -29170, -24240, -23442, -20659, -17048, -12561, -8826, 
    -3854, -654, 4204, 10249, 12725, 17381, 20918, 21801, 26591, 29079, 
    30193, 30068, 29717, 31523, 30632, 27554, 26933, 22602, 20319, 16377, 
    12209, 9001, 4444, 922, -4040, -10576, -12115, -15007, -19503, -24556, 
    -25523, -28165, -30389, -31108, -30471, -30505, -29989, -27974, -25498, 
    -23182, -20669, -15604, -12154, -8804, -4041, -1798, 4383, 9036, 11812, 
    15462, 20865, 22602, 24740, 28284, 29755, 30208, 31072, 31668, 29916, 
    28206, 25118, 23677, 20614, 17278, 12881, 8088, 5743, -500, -4846, -8264, 
    -11113, -16231, -21520, -23290, -26938, -27286, -28405, -30680, -30439, 
    -29532, -30125, -28692, -26349, -23074, -19278, -17001, -12726, -7949, 
    -3079, -860, 5262, 7097, 13222, 16790, 21376, 23300, 25592, 27748, 30353, 
    31458, 30101, 29914, 29364, 27744, 26800, 24052, 20282, 16611, 12563, 
    9197, 4730, 608, -4191, -7842, -12590, -15642, -19280, -23667, -25614, 
    -26393, -28011, -30784, -31170, -30082, -28631, -27857, -27561, -24948, 
    -19781, -16108, -12783, -10041, -5296, 882, 4112, 8378, 11176, 15814, 
    21176, 24340, 23947, 28066, 28596, 29746, 30513, 30268, 30087, 26761, 
    26206, 23089, 20412, 17653, 15037, 9180, 6191, 928, -4226, -8448, -13583, 
    -16407, -18349, -23530, -25428, -27068, -29374, -30199, -30434, -30277, 
    -28459, -28880, -26800, -24953, -21999, -18344, -13444, -10279, -6824, 
    -879, 2999, 6430, 10383, 14882, 19018, 21596, 24952, 28707, 29477, 31473, 
    30197, 30021, 30045, 29516, 28129, 24832, 20499, 18097, 13608, 8839, 
    6618, 1253, -4099, -8450, -11046, -14181, -19968, -21674, -26189, -28275, 
    -29446, -30865, -32023, -30964, -30935, -29356, -26668, -23934, -22334, 
    -18708, -14348, -11005, -4890, -1747, 3617, 8068, 11424, 15061, 18748, 
    22718, 24140, 27129, 30559, 31484, 30887, 30980, 30066, 28204, 26984, 
    24476, 23021, 18126, 15368, 9576, 5101, 1463, -2431, -6348, -9922, 
    -13331, -19173, -22143, -23435, -26521, -29301, -30019, -31475, -29586, 
    -30960, -28269, -25781, -24682, -22057, -18215, -13954, -10688, -7557, 
    -2632, 1669, 7918, 11169, 14286, 18317, 22194, 23895, 25168, 28965, 
    31363, 29866, 30830, 31622, 29519, 28142, 25457, 21965, 18329, 14419, 
    9603, 7905, 2784, -2224, -6044, -10308, -14457, -16956, -21516, -26217, 
    -26226, -28344, -30336, -31414, -30050, -30157, -27865, -27792, -23841, 
    -22514, -17518, -16137, -10898, -7062, -2885, 2125, 5267, 10537, 14720, 
    19705, 20608, 24184, 27177, 27892, 30036, 30605, 31439, 30214, 28247, 
    27967, 24934, 21975, 17080, 15151, 11293, 7275, 3742, -697, -7045, 
    -10663, -14077, -17428, -21959, -24834, -27253, -28746, -29148, -32126, 
    -31730, -31109, -30173, -27588, -25677, -20790, -18762, -13960, -12098, 
    -8040, -1654, 942, 4868, 10052, 14076, 16964, 20106, 24453, 25993, 29037, 
    29433, 31545, 31179, 29672, 28966, 28339, 26036, 22041, 19137, 14218, 
    12515, 6423, 3389, -1006, -4879, -9544, -14513, -17634, -21428, -23187, 
    -26542, -28662, -29557, -30381, -30597, -30092, -28173, -29077, -25246, 
    -23360, -18235, -14744, -11875, -7647, -3666, 1315, 5597, 8834, 13964, 
    16830, 19378, 23094, 25380, 28417, 29943, 29930, 30338, 28733, 30332, 
    29328, 26258, 22001, 18452, 17021, 11083, 7089, 4057, -1096, -5582, 
    -9794, -12878, -17335, -19900, -23035, -27985, -27646, -28689, -30430, 
    -32511, -29777, -28581, -28467, -27018, -23292, -20846, -17032, -11406, 
    -9206, -4074, 255, 4165, 8933, 12187, 16077, 19790, 24196, 25045, 27261, 
    29288, 31008, 30227, 30479, 28312, 29141, 26768, 24685, 19396, 16750, 
    12611, 8282, 3895, -560, -3778, -7647, -11941, -17585, -20290, -24281, 
    -25595, -26679, -29771, -30181, -30065, -30996, -30370, -27193, -25123, 
    -22658, -20152, -17188, -12725, -7194, -4902, -26, 4195, 7500, 12048, 
    17263, 21343, 24394, 24583, 26858, 28656, 29509, 29854, 29908, 30585, 
    27492, 25703, 22022, 18608, 15739, 12597, 10362, 4484, -206, -3964, 
    -7596, -12022, -15923, -20090, -23810, -26022, -28708, -29422, -31222, 
    -32390, -30852, -31017, -27817, -26850, -24302, -19647, -18452, -12577, 
    -7697, -4770, -679, 3417, 9864, 11744, 16792, 20073, 22531, 25030, 26810, 
    28663, 31467, 29890, 30151, 29671, 28452, 24531, 23421, 19407, 19092, 
    13028, 8925, 4353, -133, -3431, -8593, -11171, -15651, -19090, -24513, 
    -26850, -28002, -30687, -29865, -31306, -31028, -31296, -28501, -26073, 
    -24126, -19567, -17106, -14225, -8535, -6589, -1633, 3697, 7135, 12686, 
    15781, 20515, 23016, 26009, 28644, 28691, 30858, 30307, 31013, 29949, 
    29241, 28153, 23410, 20442, 16173, 13232, 9572, 5611, 1653, -2888, -8217, 
    -11649, -16154, -19769, -21493, -24538, -27201, -29370, -30073, -32107, 
    -31028, -28877, -27667, -27731, -23276, -21683, -16396, -14523, -10957, 
    -6310, -1408, 3111, 7744, 11819, 16873, 18530, 23143, 24359, 27244, 
    27692, 30443, 31436, 30642, 29531, 27955, 25033, 25159, 21366, 17985, 
    13829, 11108, 6488, 462, -2005, -7347, -11337, -15386, -20427, -21787, 
    -24806, -27649, -28037, -29666, -30398, -31615, -29907, -29136, -28061, 
    -23325, -22895, -19522, -14756, -10470, -7426, -3223, 3051, 6299, 10923, 
    14707, 20582, 21314, 23922, 27095, 28397, 31031, 30637, 30557, 28838, 
    28859, 27143, 24644, 22182, 18234, 14378, 11557, 5065, 2848, -3224, 
    -5577, -11209, -14767, -18514, -21814, -24316, -27972, -29148, -30310, 
    -30251, -29041, -29997, -28337, -26430, -25839, -21001, -17285, -14493, 
    -11457, -6804, -2174, 1265, 8316, 11822, 15072, 17801, 22816, 25418, 
    26924, 27437, 29976, 32091, 30532, 28962, 29724, 27746, 23474, 22097, 
    18089, 16376, 9834, 6391, 1297, -2452, -4919, -9653, -14861, -18318, 
    -22248, -23972, -27054, -28651, -30534, -31723, -31117, -30654, -28131, 
    -25989, -24651, -22863, -19001, -15651, -11178, -8214, -2047, 1896, 5884, 
    9183, 14693, 17908, 21796, 25544, 27200, 28279, 28917, 30845, 32658, 
    31518, 30016, 26750, 25690, 21787, 19303, 16037, 10784, 7733, 2854, 
    -1620, -6203, -8976, -13467, -19721, -21977, -25201, -25523, -27584, 
    -28919, -30554, -31022, -29013, -27934, -27032, -23872, -22005, -19733, 
    -17303, -11487, -7191, -1502, 1696, 5311, 10022, 13570, 16357, 19686, 
    23380, 25454, 28438, 29339, 29407, 29398, 30205, 28933, 26400, 26296, 
    21291, 20803, 16036, 12275, 8619, 2836, -344, -5950, -8733, -13938, 
    -17142, -20351, -24764, -27752, -28580, -29745, -29980, -32127, -29407, 
    -28858, -26695, -25318, -23293, -18579, -16824, -11595, -7482, -2146, 
    1049, 5708, 8029, 13247, 17568, 19816, 22391, 26692, 27573, 29628, 30527, 
    30034, 31047, 28741, 28452, 26527, 21301, 18608, 15383, 13160, 8733, 
    2760, 255, -5426, -9332, -12589, -16487, -21832, -23680, -26835, -27066, 
    -29666, -31682, -30557, -30190, -29638, -26868, -26113, -21492, -19907, 
    -15411, -12953, -8819, -3478, 886, 4272, 7934, 12626, 16763, 21522, 
    24199, 26101, 27311, 29398, 31459, 32181, 31337, 29888, 28892, 27239, 
    22014, 18928, 16287, 12995, 9194, 4472, -895, -4605, -10238, -13799, 
    -17554, -19767, -24959, -26997, -28170, -30146, -29140, -31260, -30451, 
    -30791, -29046, -26522, -23060, -19574, -16289, -11061, -8784, -4135, 
    -889, 5006, 8587, 13016, 16332, 19628, 21854, 26239, 28652, 29435, 29365, 
    31712, 31129, 29476, 29686, 25706, 23463, 21590, 16962, 13203, 9479, 
    3786, 86, -4393, -8685, -12576, -16407, -21454, -24049, -25639, -27227, 
    -29007, -30641, -31541, -31399, -29571, -27674, -26584, -23703, -20752, 
    -15659, -12996, -9060, -5607, 148, 3596, 6912, 13007, 16439, 20921, 
    21765, 24624, 28889, 29225, 30139, 30242, 30640, 30964, 28637, 25535, 
    25340, 20474, 17521, 13868, 9684, 5013, 969, -3531, -8591, -12563, 
    -15983, -21225, -23101, -25067, -27678, -29941, -30295, -30331, -30457, 
    -28998, -29272, -27133, -23386, -21098, -17436, -12668, -8541, -4721, 
    699, 2919, 9160, 12528, 14832, 19312, 22416, 24105, 27765, 29841, 29547, 
    30461, 31056, 30002, 28216, 26660, 24408, 20965, 17627, 13946, 10358, 
    5851, 1235, -3730, -6636, -11533, -15814, -18706, -22381, -25228, -26405, 
    -29203, -30062, -30190, -29449, -29897, -29281, -27416, -24291, -19846, 
    -19328, -13231, -8606, -6102, -1687, 4740, 8636, 12582, 15932, 19128, 
    21706, 25309, 27289, 30470, 30777, 30996, 30971, 30927, 28353, 26509, 
    25019, 19983, 17545, 12905, 9913, 7058, 1673, -3649, -7971, -12581, 
    -15833, -18142, -21905, -24755, -26793, -28041, -31176, -30045, -29659, 
    -31167, -28259, -25142, -25413, -21504, -16893, -14976, -9160, -5928, 
    -2466, 2855, 7643, 10578, 14134, 19029, 21914, 24398, 27207, 28382, 
    30437, 30488, 30088, 31644, 30391, 26524, 23885, 20520, 18693, 13844, 
    9301, 8037, 1551, -3074, -7440, -10586, -14849, -18476, -23540, -24384, 
    -26978, -28125, -29939, -30110, -31275, -30576, -29133, -28661, -25389, 
    -22520, -17785, -15373, -10980, -5339, -1923, 1037, 5884, 10715, 13561, 
    18752, 22454, 25906, 27749, 30059, 29315, 31194, 30535, 29411, 28908, 
    26518, 25460, 22354, 17897, 14454, 12348, 5817, 3055, -1735, -6269, 
    -10223, -15319, -17520, -21940, -25077, -26098, -29405, -29549, -31439, 
    -29422, -29894, -29111, -26905, -23881, -21796, -19587, -15438, -10786, 
    -6845, -3889, 3267, 5901, 10601, 14299, 19573, 19976, 23976, 28009, 
    28797, 29051, 30438, 29872, 31983, 30253, 26345, 23791, 22004, 18637, 
    15003, 11970, 7150, 1644, -581, -5915, -9498, -15024, -18579, -21242, 
    -22714, -27119, -28471, -29091, -32091, -32065, -30816, -29565, -27792, 
    -23451, -21930, -19192, -16861, -12334, -7313, -3260, 1530, 6333, 10666, 
    13680, 16468, 19601, 23942, 25766, 28470, 30278, 31011, 31145, 29361, 
    29790, 27048, 24708, 23872, 20438, 16086, 10912, 7090, 3151, -1577, 
    -6283, -9011, -14756, -16134, -21134, -22715, -26570, -29017, -28564, 
    -29586, -29810, -29416, -28902, -27206, -26078, -21259, -18819, -15732, 
    -10804, -7022, -3184, 2023, 4429, 9500, 12922, 17030, 20436, 22619, 
    26561, 27932, 30260, 29709, 31044, 29236, 29460, 27679, 24764, 23665, 
    19424, 15920, 10873, 7904, 3427, -216, -4448, -10075, -12909, -17054, 
    -20910, -22113, -26121, -27580, -28563, -29726, -32267, -28583, -29549, 
    -26995, -26275, -21905, -18875, -16202, -12626, -7498, -3566, 328, 3897, 
    10379, 13564, 17116, 20004, 23046, 25056, 28268, 29776, 28701, 30927, 
    29725, 29601, 27418, 24663, 22438, 20067, 14906, 12850, 8322, 4461, 96, 
    -5500, -7458, -12192, -17539, -20128, -25139, -25220, -28874, -30438, 
    -30580, -31049, -31516, -29847, -28229, -26089, -22795, -19106, -17394, 
    -13070, -7934, -5595, 786, 4773, 7840, 13396, 14907, 20170, 23540, 24793, 
    27878, 29791, 30877, 31777, 30505, 29994, 27244, 24735, 22679, 21158, 
    15836, 13056, 7876, 4749, -1552, -2796, -7906, -11308, -15565, -19742, 
    -22381, -25877, -26651, -29192, -30321, -31276, -31788, -30046, -28802, 
    -27237, -22847, -22158, -16380, -13179, -9842, -5126, 440, 4479, 8789, 
    11659, 16687, 20883, 23706, 24428, 26814, 29587, 28856, 30650, 29846, 
    30428, 27212, 27669, 23863, 20756, 17762, 13951, 8796, 4702, 508, -3389, 
    -6364, -12636, -16030, -19846, -20962, -26268, -27798, -30137, -29690, 
    -31094, -31151, -29088, -27384, -25692, -24672, -22086, -17445, -11893, 
    -8601, -5953, -2288, 4194, 6450, 11777, 16869, 19295, 22203, 24844, 
    26733, 28308, 30466, 30206, 30890, 30766, 27129, 25243, 23409, 20630, 
    17175, 13375, 9645, 3808, 733, -3418, -7422, -10995, -15014, -19835, 
    -22700, -24548, -28324, -29179, -31072, -30831, -30580, -29617, -29767, 
    -26189, -25134, -20555, -16589, -14271, -10745, -4432, -1308, 3131, 6317, 
    10017, 16424, 20027, 21816, 24124, 26478, 29876, 31232, 32248, 31884, 
    30550, 28711, 25348, 22926, 20493, 18405, 14587, 10134, 5082, 1042, 
    -2854, -6387, -10081, -15605, -19061, -22228, -25095, -26771, -28498, 
    -30292, -30976, -31524, -29890, -28509, -26099, -23915, -22149, -17613, 
    -14855, -10935, -5685, -2346, 3923, 6916, 10888, 15540, 19712, 22348, 
    23708, 26883, 28020, 31100, 30737, 31470, 30038, 29445, 28031, 24295, 
    23449, 18257, 14432, 9617, 5427, 1769, -1288, -5867, -10237, -15077, 
    -17975, -21124, -23854, -26455, -29445, -30249, -30645, -29900, -29779, 
    -29702, -27031, -24753, -20443, -17577, -14631, -10224, -5302, -2103, 
    3978, 7290, 10906, 15521, 18227, 22775, 24340, 27339, 29669, 31236, 
    29609, 29633, 28824, 27661, 28227, 23301, 21469, 19352, 14355, 10938, 
    6888, 1877, -1988, -5604, -10337, -13920, -17800, -21154, -25264, -26513, 
    -27847, -29799, -30424, -29973, -29478, -29701, -27460, -25546, -21495, 
    -18030, -15114, -11484, -6505, -2880, 1867, 6227, 9148, 14376, 17818, 
    22884, 23454, 27685, 29276, 30326, 30947, 30062, 29802, 29035, 27757, 
    24164, 21229, 19608, 15379, 12117, 6023, 2539, -2832, -6415, -10128, 
    -13699, -16821, -19946, -24702, -27046, -29238, -30590, -29864, -29579, 
    -30635, -29250, -27507, -24464, -21181, -19220, -16802, -11433, -6728, 
    -4344, 1274, 4882, 9496, 15508, 17812, 20574, 23776, 27681, 29300, 30130, 
    30431, 32345, 30986, 29301, 29311, 24432, 22806, 18776, 16467, 11171, 
    8091, 2492, -1338, -4875, -9179, -13461, -16854, -20747, -24424, -26991, 
    -27640, -30807, -31276, -31110, -30213, -28674, -28387, -24606, -21876, 
    -18684, -16199, -10655, -7974, -3597, 882, 5039, 8819, 14555, 18595, 
    20307, 23915, 27924, 27163, 30810, 29822, 31428, 30434, 27567, 28033, 
    24653, 23154, 18620, 14367, 12379, 7674, 2598, -178, -4073, -10221, 
    -14392, -16637, -21306, -24761, -26339, -27607, -31044, -30457, -29653, 
    -30371, -29387, -28432, -25552, -24362, -20039, -16915, -12405, -8237, 
    -5414, 1248, 4926, 7973, 12956, 17309, 21633, 24018, 26417, 28936, 29681, 
    31434, 30217, 30709, 29424, 27872, 25901, 22981, 20696, 16560, 12642, 
    7716, 4094, 440, -3445, -9335, -11358, -17304, -20706, -23541, -26930, 
    -27854, -28986, -29209, -30770, -29397, -28098, -29350, -25097, -24110, 
    -20875, -15966, -12233, -8964, -3823, -464, 4274, 8727, 13513, 16665, 
    18919, 23192, 24335, 27541, 29170, 30206, 30281, 31175, 28194, 28297, 
    24876, 23429, 19748, 16794, 12592, 8902, 6374, 162, -2703, -8042, -12144, 
    -16755, -18942, -23799, -25913, -26790, -30174, -30920, -29898, -30621, 
    -29011, -27383, -27330, -23596, -20587, -15882, -13328, -9385, -4992, 
    -702, 3070, 8241, 11623, 17754, 19994, 22234, 25516, 27129, 28762, 30524, 
    31819, 29528, 28457, 28017, 27933, 24198, 19930, 16791, 13655, 8279, 
    4257, 1258, -4314, -8353, -12479, -16123, -18894, -22525, -25285, -26559, 
    -30052, -30749, -31092, -30441, -31229, -28309, -25899, -23712, -20898, 
    -15839, -13187, -9111, -3948, 358, 3668, 6684, 13194, 16207, 19636, 
    22018, 23761, 28093, 30061, 31497, 31184, 30623, 28258, 28202, 27736, 
    23145, 21406, 16355, 12648, 9042, 6177, 1135, -2855, -6383, -12364, 
    -15087, -19087, -23208, -24397, -27861, -29561, -31602, -29343, -30141, 
    -28326, -27922, -26667, -23462, -21043, -18906, -14133, -11224, -6496, 
    -2074, 2760, 6574, 13228, 15414, 19196, 21382, 26610, 27135, 29682, 
    29206, 31525, 29545, 30008, 29430, 26027, 25098, 22001, 18557, 13396, 
    10425, 5207, 1913, -4009, -7824, -11481, -15438, -18606, -21689, -24622, 
    -27209, -29859, -31408, -30299, -30721, -29760, -27998, -26116, -24004, 
    -21224, -18356, -12886, -10280, -6896, -1317, 2241, 7759, 10837, 15895, 
    18541, 20361, 24196, 26585, 29179, 30143, 29619, 31104, 29496, 28084, 
    26801, 22990, 20321, 18862, 14537, 10668, 6000, 1987, -1292, -6973, 
    -10963, -13472, -18589, -21616, -24776, -28274, -27482, -30341, -29660, 
    -32092, -30313, -27462, -27204, -25424, -20705, -17500, -13994, -11932, 
    -6879, -2445, 2124, 5776, 12104, 13923, 19161, 20992, 25644, 27669, 
    28925, 29191, 29440, 31969, 31636, 29821, 27006, 23196, 22257, 19080, 
    14345, 11490, 6512, 2664, -1840, -5126, -9783, -16196, -18387, -21263, 
    -24817, -26496, -27523, -30744, -29988, -30811, -28599, -29611, -26525, 
    -25920, -22232, -18939, -16504, -10242, -5963, -1334, 2686, 7258, 11105, 
    13271, 19029, 21796, 25003, 27186, 29279, 29845, 29956, 31387, 30751, 
    29458, 28177, 25684, 21751, 19394, 16989, 10369, 6458, 2660, -227, -6121, 
    -9422, -13302, -16102, -22189, -24184, -27231, -28135, -29752, -30800, 
    -29965, -28573, -28427, -27222, -25389, -21396, -18156, -16682, -12152, 
    -7817, -3026, 282, 3989, 11228, 13118, 16674, 21511, 25021, 25352, 27382, 
    28997, 29950, 29840, 31166, 29288, 28120, 25072, 21893, 19678, 16944, 
    11805, 7519, 3743, -1339, -4603, -9285, -13787, -17364, -20908, -24512, 
    -27460, -26876, -29927, -30775, -32050, -29843, -28426, -27150, -25572, 
    -23675, -20942, -17049, -11905, -7672, -3703, 2129, 4827, 9097, 13008, 
    18685, 20377, 25435, 25399, 29017, 28429, 30396, 31042, 30410, 29669, 
    27669, 26735, 22474, 20282, 15960, 12825, 7212, 4276, -992, -3930, 
    -10410, -15026, -17420, -22417, -23129, -25181, -27568, -30904, -32447, 
    -32342, -32111, -30001, -26914, -24894, -23105, -18535, -16467, -12570, 
    -7436, -4203, 1718, 4909, 9105, 13397, 17535, 18991, 22434, 24901, 28880, 
    30265, 30533, 29881, 31063, 28864, 29189, 25492, 22620, 20416, 16194, 
    13246, 9791, 3881, -63, -3463, -7964, -13127, -16705, -21169, -24506, 
    -25413, -28198, -29320, -31781, -30227, -30339, -30813, -28724, -25423, 
    -22246, -19615, -16252, -13114, -9895, -4590, 394, 4927, 8309, 13786, 
    15602, 20578, 23196, 26046, 27308, 30006, 31223, 30947, 30762, 30158, 
    28752, 26597, 22933, 19929, 16784, 13820, 9412, 5727, 319, -3830, -9528, 
    -11853, -15562, -19467, -23065, -25290, -26782, -28952, -29649, -31326, 
    -29868, -31533, -27915, -26729, -23480, -20590, -17074, -13418, -9547, 
    -5070, 1231, 4659, 9976, 12328, 15652, 21101, 23003, 26011, 27064, 30457, 
    31976, 31615, 31138, 29060, 29211, 25378, 23252, 20593, 17677, 13877, 
    7861, 4684, 1169, -4911, -9124, -12594, -15246, -21060, -23389, -26875, 
    -27743, -29936, -30170, -30644, -30917, -30427, -28312, -26039, -22749, 
    -19119, -16310, -13945, -11089, -5413, -1458, 3734, 7523, 12676, 16649, 
    18328, 22691, 24312, 27711, 27953, 31408, 31822, 30722, 29168, 27520, 
    25323, 23832, 21081, 17166, 14319, 8394, 6116, 1694, -2360, -6482, 
    -10631, -15546, -19414, -23978, -25165, -27362, -28210, -29819, -31209, 
    -31050, -30092, -28916, -26674, -25132, -20357, -17586, -13993, -11502, 
    -6824, -54, 3944, 8748, 12912, 16874, 18463, 22280, 23852, 27264, 29195, 
    29131, 29786, 30986, 30344, 28783, 26463, 24080, 21168, 18631, 14289, 
    9165, 5299, 721, -4047, -7302, -11346, -14837, -19498, -22893, -23826, 
    -26959, -29049, -30366, -30140, -30081, -31043, -30493, -25584, -24019, 
    -22310, -19391, -14260, -11751, -6533, -2592, 1259, 7128, 11438, 14614, 
    17044, 21909, 23723, 27246, 28735, 29102, 30818, 30199, 30006, 28710, 
    26934, 22749, 21576, 17386, 13187, 9721, 5234, 1500, -2292, -6551, -9986, 
    -16425, -17307, -21931, -24160, -27102, -29980, -28934, -30485, -31591, 
    -29715, -29076, -26624, -25426, -21083, -17796, -14120, -11482, -6449, 
    -1953, 2699, 7033, 10457, 14186, 18187, 20330, 25092, 27542, 28728, 
    30842, 30397, 30462, 29751, 28645, 25945, 25428, 21365, 18124, 14168, 
    11204, 6769, 2435, -2936, -5266, -10762, -14031, -18727, -21563, -24324, 
    -28133, -27502, -29973, -30204, -31295, -30521, -27424, -27129, -26200, 
    -22488, -19383, -15179, -11994, -6779, -1904, 1856, 5708, 9248, 13982, 
    18412, 22630, 24981, 26598, 27111, 31821, 29792, 30584, 29863, 28704, 
    26303, 24326, 22626, 18836, 15444, 12177, 7934, 2863, -487, -4534, -9551, 
    -14666, -18084, -20258, -24822, -27302, -30141, -30472, -31092, -31185, 
    -31201, -29475, -26326, -25711, -23005, -19659, -15610, -11897, -7886, 
    -2806, 2529, 5856, 10555, 13479, 19082, 22220, 23123, 26957, 28601, 
    29343, 29821, 32125, 31074, 28226, 26698, 26175, 21092, 19509, 16697, 
    11739, 6704, 4470, -396, -3825, -10070, -13416, -17991, -22054, -24799, 
    -28051, -29210, -30941, -30667, -30828, -30038, -29466, -26487, -24439, 
    -22348, -20843, -16641, -11057, -8774, -3364, -855, 4422, 9009, 13908, 
    17029, 21188, 24491, 26721, 29957, 29741, 31897, 31338, 30034, 29611, 
    27135, 25209, 23455, 20625, 17203, 12140, 9074, 4442, 937, -5662, -9488, 
    -13403, -16633, -19356, -22690, -26443, -28379, -29387, -30140, -30819, 
    -31612, -28737, -28715, -26946, -22888, -20975, -15928, -11121, -7958, 
    -4809, 1346, 4205, 10141, 12642, 17974, 19078, 23808, 26053, 28071, 
    29876, 30824, 30047, 29816, 30014, 28032, 26202, 23387, 21175, 17366, 
    11225, 7535, 3675, -1242, -5219, -7808, -13199, -14990, -20922, -23182, 
    -25307, -27072, -29368, -31153, -30876, -31661, -29707, -29231, -25877, 
    -23767, -21012, -16929, -12648, -8750, -3880, -165, 5548, 8122, 12602, 
    16447, 20622, 24578, 25435, 29527, 29218, 30410, 32445, 30544, 30045, 
    28843, 26198, 23736, 20063, 15878, 13786, 9546, 4794, 909, -3723, -8051, 
    -12219, -16747, -20084, -21356, -25532, -27690, -29117, -31101, -30378, 
    -31577, -30326, -29730, -27279, -23235, -20740, -15500, -12732, -9464, 
    -5769, -2234, 5337, 7689, 13727, 16028, 19660, 22645, 27330, 28550, 
    29818, 31402, 29745, 29207, 30325, 30074, 26864, 23226, 20930, 18060, 
    13304, 9221, 5783, -244, -2920, -7172, -10763, -15115, -19809, -22291, 
    -25634, -27753, -30565, -30592, -31316, -32026, -30684, -28822, -25856, 
    -23441, -21002, -16061, -12803, -9651, -6409, -1069, 3248, 6741, 11698, 
    16050, 19501, 22302, 25678, 27269, 29939, 30591, 30987, 30668, 29490, 
    28981, 24960, 24076, 20923, 18438, 14020, 10933, 4809, 1860, -3899, 
    -6932, -10555, -15092, -19392, -22270, -23733, -28080, -29433, -31653, 
    -30084, -30914, -30390, -29469, -25439, -24040, -20594, -17218, -15302, 
    -10997, -6384, -2608, 1724, 7581, 11752, 15338, 19753, 22754, 24084, 
    26306, 28876, 31090, 31168, 30989, 29503, 28410, 25658, 25509, 22312, 
    17839, 13624, 9744, 6478, 2819, -4467, -7743, -9916, -15417, -19109, 
    -21590, -23933, -27868, -29123, -30628, -31137, -31577, -30302, -29450, 
    -26864, -24057, -21410, -17249, -14945, -8993, -5867, -2285, 1542, 6318, 
    10903, 13481, 18234, 21609, 24341, 28491, 27376, 28802, 31357, 31335, 
    28793, 27616, 26225, 24560, 20311, 18582, 12694, 10164, 6249, 455, -2844, 
    -6893, -11111, -14322, -19546, -20355, -25654, -28005, -29835, -30965, 
    -30017, -30078, -30890, -27832, -26089, -24242, -22405, -20122, -13863, 
    -10340, -5874, -2208, 2744, 5065, 10758, 13590, 18200, 21746, 24212, 
    26557, 27623, 29509, 31128, 30060, 30472, 28192, 28358, 24168, 21476, 
    19242, 13922, 11422, 5459, 3628, -1831, -5019, -10668, -13833, -17500, 
    -20579, -25162, -27118, -29818, -29300, -29923, -32128, -31054, -28057, 
    -26380, -24084, -21839, -18643, -15793, -11989, -8078, -1595, 3137, 6207, 
    10441, 14846, 17623, 22158, 24416, 27272, 28796, 30475, 32147, 31738, 
    30637, 27814, 28676, 25234, 20833, 18584, 15020, 11661, 6405, 3656, 
    -1810, -7269, -9636, -12882, -17940, -21019, -23367, -25849, -29076, 
    -29220, -31563, -31637, -29389, -27909, -27667, -25124, -21935, -18921, 
    -14961, -11749, -7318, -3270, 2129, 6145, 10669, 14265, 17392, 19982, 
    25430, 26474, 28006, 28790, 31571, 30510, 29491, 29067, 28135, 24026, 
    23216, 19063, 14749, 11668, 6958, 3534, -2016, -5464, -10705, -12587, 
    -17281, -22195, -24422, -25835, -27690, -28324, -31240, -30554, -31764, 
    -29392, -28055, -25065, -24307, -20619, -14588, -11616, -7918, -5075, 
    2143, 6079, 9582, 13828, 17395, 21746, 23806, 26412, 28499, 29215, 30506, 
    29813, 30330, 28350, 27375, 26592, 23291, 20080, 16519, 12273, 8297, 
    3929, -325, -5496, -10002, -14228, -18255, -20236, -25079, -27184, 
    -28557, -29068, -31116, -31997, -32172, -29672, -27742, -25943, -21981, 
    -20995, -14791, -13807, -7460, -3450, -171, 4774, 7795, 13512, 17919, 
    21080, 23532, 25368, 27969, 28233, 30324, 30566, 30260, 29548, 27403, 
    25742, 23978, 20497, 15949, 13212, 8543, 4218, 620, -4647, -8780, -11882, 
    -16108, -20666, -23957, -26466, -28922, -30673, -30495, -29960, -30997, 
    -29987, -27626, -25306, -24966, -21400, -16510, -11454, -8249, -3297, 
    101, 4481, 9081, 13544, 16692, 20681, 23604, 24292, 27726, 28682, 30416, 
    30510, 29875, 30026, 27849, 26171, 23287, 20655, 17106, 13440, 9507, 
    4999, 405, -4394, -8151, -12750, -16379, -19605, -23544, -24884, -27956, 
    -29305, -31234, -30635, -30441, -29492, -28358, -27329, -24088, -20638, 
    -16214, -12827, -7880, -5056, 552, 2757, 8909, 12306, 15169, 18768, 
    24539, 27130, 27798, 30622, 31316, 30844, 30781, 29448, 28613, 26290, 
    23989, 21964, 17144, 12909, 9379, 6225, -400, -4252, -8121, -11343, 
    -14291, -20467, -22946, -25297, -27050, -28428, -29995, -31426, -30447, 
    -29321, -27973, -27161, -25301, -20469, -16629, -13551, -9729, -5821, 
    -1307, 3206, 7765, 11490, 16511, 20334, 22736, 25091, 27376, 29454, 
    29557, 30718, 30690, 28386, 29094, 24878, 25309, 22116, 17690, 13873, 
    10430, 4846, -66, -1953, -7180, -10770, -17403, -18089, -22793, -23873, 
    -28630, -30231, -30449, -31573, -30925, -29355, -27762, -26914, -24205, 
    -21903, -16593, -14033, -10618, -6798, -1295, 2469, 8421, 11094, 15368, 
    18763, 21858, 25167, 26707, 31056, 29512, 30948, 31641, 30361, 28880, 
    27224, 23860, 21481, 18226, 13896, 10728, 5576, 2080, -1865, -6220, 
    -9548, -16247, -18332, -22857, -25572, -27726, -29490, -30685, -29634, 
    -30577, -29350, -28916, -26820, -23852, -21959, -18862, -14035, -10320, 
    -5715, -1715, 1934, 6920, 9731, 16278, 17778, 22335, 25656, 28501, 29520, 
    29522, 31421, 30217, 29747, 27939, 27466, 25735, 21241, 16775, 13963, 
    10877, 7849, 2930, -2527, -7122, -10280, -15715, -17361, -22098, -25110, 
    -27295, -29265, -28601, -31200, -30120, -30566, -29653, -26621, -23835, 
    -22569, -17039, -13570, -9920, -5227, -1688, 1509, 6353, 12234, 14679, 
    19830, 22045, 24267, 27206, 29081, 30827, 29960, 30648, 30324, 30216, 
    27381, 25088, 22977, 17886, 14409, 10589, 5898, 2111, -2163, -6011, 
    -9361, -14462, -18321, -21129, -25354, -26870, -27958, -29726, -29863, 
    -32066, -30114, -28673, -27440, -25453, -22504, -17986, -14292, -10632, 
    -6298, -3519, 674, 6879, 9573, 14356, 17946, 20403, 23775, 26939, 28655, 
    30476, 30411, 30162, 30298, 29254, 27471, 24974, 21944, 18719, 16234, 
    10561, 7778, 4127, -787, -6409, -10521, -15878, -19375, -21310, -23154, 
    -27205, -28232, -30251, -31428, -31310, -31308, -29079, -26348, -23733, 
    -23357, -18034, -15521, -11183, -7870, -2044, 968, 6872, 10752, 15244, 
    18132, 20010, 23594, 25883, 29193, 29300, 28871, 31103, 30132, 28324, 
    27273, 24684, 23180, 18008, 16053, 11963, 7262, 4461, -865, -5677, -9674, 
    -14280, -17734, -20401, -22866, -27663, -28901, -29718, -30031, -31440, 
    -31211, -29202, -28932, -25205, -22430, -20546, -16603, -11496, -7039, 
    -3630, 252, 5570, 10094, 12411, 16625, 22004, 22535, 25487, 28907, 29681, 
    30533, 31164, 30210, 28943, 29089, 26005, 24091, 18669, 16144, 13465, 
    7723, 4356, -672, -5270, -9434, -14653, -18107, -20386, -23170, -26004, 
    -29003, -28634, -29454, -30461, -30037, -29445, -27356, -27305, -23580, 
    -18940, -15865, -12980, -7473, -4848, 67, 5190, 8443, 13999, 17456, 
    20896, 22998, 25547, 27709, 28949, 29111, 30624, 29930, 30600, 27607, 
    25401, 21814, 18302, 14559, 11685, 8608, 3715, 194, -5919, -8814, -13973, 
    -16335, -20243, -23779, -24517, -28435, -28506, -31855, -30304, -31308, 
    -27951, -27485, -25464, -23309, -21038, -15873, -13476, -8901, -4648, 
    -1095, 4830, 8634, 12009, 16486, 20327, 23048, 26594, 27299, 29774, 
    30475, 29390, 30216, 29976, 28208, 25151, 23986, 20542, 18086, 12793, 
    8910, 5197, 638, -5251, -9006, -12192, -16563, -20835, -22948, -24955, 
    -27165, -30449, -30904, -31295, -30845, -30371, -27923, -26514, -22582, 
    -19464, -17546, -14347, -8723, -5399, -1397, 3576, 8518, 12886, 16079, 
    21118, 23514, 24033, 28801, 28712, 29166, 29392, 29703, 29400, 27841, 
    26488, 24032, 20694, 17771, 12558, 10170, 4198, 1325, -3656, -7934, 
    -12037, -15868, -18640, -23226, -23971, -26843, -28406, -30651, -30972, 
    -31528, -29018, -28676, -25655, -23597, -20854, -16648, -14443, -9967, 
    -4654, -1411, 5064, 7112, 11218, 15915, 18545, 22985, 27025, 27989, 
    29522, 31067, 30630, 30161, 29276, 28460, 26168, 24572, 20017, 18405, 
    12815, 9253, 5583, -377, -2890, -7008, -11529, -16563, -19407, -22141, 
    -24574, -27092, -28160, -29901, -31194, -31297, -31088, -28658, -26663, 
    -25093, -21109, -16375, -14294, -10270, -4927, -638, 2143, 6377, 11561, 
    15039, 18572, 23943, 24440, 27501, 28775, 30882, 30660, 29768, 31677, 
    28607, 28068, 23408, 22029, 18915, 14133, 10087, 6860, 1599, -3190, 
    -8595, -12530, -15688, -19247, -20882, -24764, -28092, -27940, -30398, 
    -30148, -31102, -29072, -29495, -27606, -23972, -21975, -17064, -12977, 
    -10793, -6442, -2294, 1838, 6679, 10915, 15318, 18629, 22892, 24171, 
    27200, 30150, 29945, 29393, 31437, 29859, 28092, 25181, 26217, 22512, 
    17540, 13824, 9657, 6170, 480, -2846, -6237, -12281, -16333, -17321, 
    -21779, -24134, -25902, -28664, -29954, -30429, -31668, -29954, -28155, 
    -28418, -25190, -20867, -18048, -13272, -12018, -6213, -1089, 1264, 7589, 
    9831, 14725, 18957, 21354, 25872, 27657, 29088, 30231, 31497, 31249, 
    30315, 30263, 27734, 23807, 22333, 18472, 15129, 10705, 7813, 3193, 
    -2124, -6437, -10984, -14219, -19269, -22409, -25129, -25740, -27191, 
    -31595, -30093, -30748, -30473, -27577, -27298, -24906, -20646, -18092, 
    -15642, -11970, -7318, -2585, 1914, 6263, 9461, 13729, 17968, 20848, 
    24318, 27306, 28042, 29808, 30784, 29684, 31605, 30171, 28662, 23283, 
    22297, 18560, 14551, 12574, 7881, 2033, 84, -6239, -10149, -13885, 
    -17842, -21830, -23133, -26592, -27536, -29881, -31682, -30576, -31746, 
    -28319, -27318, -25246, -22375, -20150, -14621, -10750, -7282, -2221, 
    2072, 5047, 10065, 15370, 18752, 21274, 23935, 26897, 27936, 29476, 
    31071, 30739, 29885, 29474, 28814, 24314, 23353, 18822, 15875, 11294, 
    8535, 4123, -583, -6257, -9471, -14290, -16735, -21482, -24246, -27715, 
    -29256, -28818, -32322, -30255, -29111, -30436, -27966, -24242, -22447, 
    -19167, -15140, -11693, -6388, -3714, 421, 4994, 8998, 15127, 17614, 
    20730, 23692, 27617, 28841, 29192, 31547, 30824, 31750, 29466, 28655, 
    26017, 22408, 19883, 16548, 10819, 8496, 4042, 80, -4782, -10047, -14316, 
    -16072, -20728, -24686, -25872, -27985, -29137, -31780, -30311, -29670, 
    -29999, -26895, -25734, -23800, -19464, -16308, -13249, -8689, -4879, 
    1097, 4726, 7979, 13641, 17385, 20699, 22884, 26813, 28236, 29858, 31114, 
    30503, 31579, 29440, 27246, 25561, 23219, 18913, 16836, 12428, 8585, 
    4553, 1203, -4017, -10280, -12942, -15844, -18733, -23703, -26681, 
    -28099, -29682, -31287, -29931, -29486, -29713, -27976, -26411, -24310, 
    -21577, -17027, -13060, -9904, -3388, 769, 4637, 10111, 11426, 16938, 
    21024, 24493, 24847, 28491, 30716, 30274, 30188, 29246, 28480, 28519, 
    26035, 23473, 19646, 16889, 11386, 8991, 5738, 196, -5139, -8121, -13775, 
    -17903, -18759, -23385, -27294, -28694, -31228, -30929, -30538, -30157, 
    -30568, -28477, -26673, -23148, -21184, -16292, -14432, -9136, -4961, 
    -1450, 2849, 6725, 10910, 15757, 20223, 22500, 25681, 28315, 30153, 
    28652, 31193, 31753, 30638, 27618, 26310, 24696, 20566, 17165, 12576, 
    9974, 5332, 1450, -1912, -7661, -12594, -16767, -19334, -23121, -26759, 
    -27499, -29095, -29430, -30127, -30602, -29834, -28091, -26414, -23748, 
    -20218, -17843, -13864, -9391, -4815, -412, 2311, 6486, 12117, 14126, 
    19215, 21774, 25271, 27333, 29919, 29824, 32408, 31091, 30173, 27869, 
    25980, 24198, 20077, 18388, 14540, 10106, 6317, 1222, -3931, -6805, 
    -12577, -14256, -19533, -22305, -25219, -27242, -29615, -30282, -31686, 
    -30990, -29245, -28747, -25208, -23636, -20949, -17836, -14351, -10833, 
    -4601, -1230, 3858, 7652, 11785, 14796, 20652, 22466, 26718, 28222, 
    29111, 30081, 30375, 30184, 29385, 28101, 27851, 24014, 21192, 19077, 
    14418, 11820, 6555, 3142, -2053, -8718, -10851, -15156, -18893, -21612, 
    -25541, -26960, -30126, -30861, -30742, -31325, -30050, -29056, -26823, 
    -24208, -22527, -18238, -13875, -10329, -6502, -3074, 2617, 6774, 9762, 
    14427, 20029, 23371, 23822, 26706, 29355, 30049, 30541, 29484, 30654, 
    28901, 26380, 25749, 22148, 18409, 14325, 10912, 7365, 2135, -2324, 
    -6574, -10827, -13658, -19772, -20848, -23760, -27372, -30553, -29515, 
    -30577, -30532, -30521, -28986, -26783, -25417, -21851, -19337, -15775, 
    -11227, -7797, -2845, 3408, 6911, 11008, 13991, 17645, 22852, 24966, 
    28271, 29797, 30279, 30812, 30564, 31916, 28711, 26683, 24957, 22053, 
    18613, 13673, 10835, 6079, 2835, -2102, -7653, -9721, -15269, -18524, 
    -21183, -25279, -27058, -29937, -29239, -30743, -29888, -29764, -29166, 
    -27573, -24858, -20799, -18592, -16299, -12215, -7603, -1307, 649, 5920, 
    9648, 15093, 16503, 21226, 24033, 25535, 29344, 30215, 31828, 31463, 
    29400, 29094, 28098, 24448, 22186, 19081, 16521, 11230, 7518, 2539, 
    -1634, -5447, -9895, -12569, -16600, -22040, -24639, -26857, -29276, 
    -30220, -29657, -31139, -30059, -28753, -27160, -27041, -22268, -19647, 
    -15922, -10292, -6306, -1899, 2472, 5650, 11406, 13833, 17760, 20713, 
    25267, 27587, 28452, 28649, 29273, 29315, 29613, 27911, 26688, 25743, 
    22911, 19734, 15135, 11528, 7803, 2823, -2539, -4726, -11256, -13923, 
    -18529, -22358, -24619, -27011, -29011, -30578, -29621, -29240, -29997, 
    -29601, -27416, -25942, -22796, -18541, -15641, -11979, -7432, -4241, 
    -36, 7031, 8883, 13649, 15717, 21031, 22948, 26664, 28472, 29489, 30950, 
    32191, 29737, 29465, 26976, 25873, 22059, 20000, 15821, 12116, 6823, 
    5112, -911, -4335, -8021, -14363, -16776, -20383, -22817, -26720, -28960, 
    -29597, -30682, -30885, -31687, -29273, -29426, -26917, -23185, -19537, 
    -15685, -13934, -8334, -3927, 1972, 4683, 8856, 14340, 15612, 20300, 
    23318, 24587, 28560, 29590, 30625, 29684, 30580, 28917, 27936, 27287, 
    22525, 19256, 17610, 11141, 8545, 3845, -372, -3809, -9285, -13630, 
    -17911, -19806, -23946, -26134, -28716, -31396, -30792, -30723, -30961, 
    -30067, -27338, -26338, -24047, -18417, -16644, -13201, -8865, -4468, 
    -529, 4368, 8541, 12253, 15971, 19391, 23293, 27608, 27956, 31315, 31906, 
    29036, 31551, 31181, 27926, 25909, 23846, 20667, 17689, 12469, 9186, 
    4401, 1605, -4616, -9558, -11334, -16774, -18857, -21549, -26876, -26615, 
    -29683, -30349, -30860, -29443, -29095, -27966, -26707, -23789, -19276, 
    -17221, -12119, -8874, -4483, -599, 4965, 8302, 11674, 15737, 19925, 
    21699, 27184, 27740, 29385, 30831, 30575, 30981, 30480, 27188, 25910, 
    23010, 20942, 18277, 11798, 8235, 5564, 1644, -4143, -6418, -10431, 
    -15835, -19353, -22948, -25300, -28878, -29893, -29450, -31656, -31565, 
    -30246, -28118, -25029, -24854, -20727, -18262, -13980, -8130, -6706, 
    -268, 3272, 6384, 10420, 16993, 19858, 22281, 24939, 28251, 30279, 31005, 
    31781, 29834, 30212, 27930, 26783, 24481, 20971, 17467, 13385, 9240, 
    4825, 1208, -1809, -6995, -11420, -15892, -20663, -22187, -25635, -28164, 
    -29087, -31460, -30804, -30396, -29402, -29343, -25018, -24893, -20075, 
    -17611, -13379, -10619, -4204, -993, 4191, 8701, 10273, 15591, 18293, 
    22587, 24123, 27941, 30301, 31042, 28962, 31069, 31250, 28083, 27430, 
    24502, 20439, 19024, 13222, 8477, 7068, 1339, -1784, -5792, -10928, 
    -15022, -19998, -22086, -24505, -27296, -29346, -29573, -30665, -30884, 
    -31252, -27893, -26441, -23983, -19930, -17053, -14215, -9882, -5924, 
    -2368, 3157, 7058, 11323, 16515, 19811, 21829, 24473, 27585, 28176, 
    30957, 30063, 30710, 31411, 28180, 25880, 25968, 21669, 18359, 14783, 
    10325, 5595, 2741, -2589, -5734, -12457, -15784, -17076, -21750, -23104, 
    -26563, -28344, -28842, -30543, -30839, -29659, -28500, -28572, -24550, 
    -21674, -18115, -15171, -9851, -6371, -3256, 1179, 7392, 9746, 15745, 
    16924, 22412, 26281, 26218, 29391, 30303, 30104, 31789, 30265, 29977, 
    26271, 23701, 21312, 19145, 15146, 11072, 5392, 3412, -785, -6689, 
    -10386, -15441, -19258, -20157, -24333, -25089, -27902, -29832, -31093, 
    -31547, -31265, -29468, -26350, -24001, -21396, -20303, -15109, -11154, 
    -6306, -1480, 1872, 7029, 10633, 14666, 16771, 21264, 24286, 28276, 
    28634, 29696, 30798, 30554, 29576, 28745, 25953, 24192, 22938, 18307, 
    15865, 11372, 7046, 3598, -974, -6112, -9463, -14129, -18051, -20204, 
    -24590, -26596, -27473, -30234, -29523, -31365, -31009, -29653, -26453, 
    -25344, -21833, -19783, -16988, -11525, -6711, -3696, 2175, 4467, 9235, 
    14552, 18698, 22060, 22446, 26882, 28720, 29929, 30547, 31378, 31318, 
    28417, 27325, 24067, 23870, 19720, 15882, 12681, 7683, 2449, -1040, 
    -6010, -9771, -13818, -16575, -21584, -23527, -26206, -27825, -28933, 
    -30793, -31487, -30871, -30082, -26945, -26904, -21487, -20273, -16754, 
    -10599, -7151, -4677, 2030, 4797, 8658, 12514, 16667, 19755, 24902, 
    27508, 27897, 28640, 31444, 32013, 31310, 29035, 27840, 24969, 22913, 
    18247, 15618, 11267, 7224, 3939, -1166, -4859, -9704, -11921, -18705, 
    -19987, -24576, -24942, -29394, -30537, -32142, -30526, -31900, -30244, 
    -28491, -26133, -21705, -19087, -17944, -13220, -8466, -4001, 1906, 3261, 
    9848, 12512, 18626, 21536, 24514, 24477, 28068, 30109, 30245, 31677, 
    29853, 29243, 27002, 26596, 21764, 18271, 16674, 13091, 10297, 4781, 
    -1701, -3599, -9408, -12871, -16707, -20379, -24321, -25281, -29164, 
    -30971, -29421, -29282, -30628, -30672, -28576, -25858, -24554, -20928, 
    -15701, -11889, -8227, -5717, -164, 5255, 8885, 12542, 16826, 20683, 
    23952, 27524, 28914, 29292, 30215, 30899, 30239, 30257, 27051, 25081, 
    24000, 20663, 17180, 13242, 8205, 5208, 432, -4338, -8883, -12989, 
    -16318, -19686, -23705, -25243, -27766, -28823, -29788, -30200, -29544, 
    -30197, -27860, -25451, -23381, -21039, -18215, -14374, -8292, -2987, 
    -373, 5012, 9316, 12752, 15980, 18490, 23263, 25665, 27356, 30375, 31129, 
    30848, 30926, 29627, 27329, 26415, 23851, 18959, 16357, 13744, 10950, 
    5639, 1264, -3719, -8512, -11098, -15648, -19097, -22251, -26583, -27330, 
    -29387, -29884, -31445, -30591, -29525, -27316, -26098, -23028, -19952, 
    -18073, -13508, -9274, -3983, -840, 2695, 6811, 11366, 16177, 18524, 
    22493, 24455, 26268, 29835, 30444, 30271, 30829, 30051, 27868, 26380, 
    23649, 20342, 16664, 13680, 10751, 6759, 156, -4266, -6200, -11846, 
    -15674, -19386, -22480, -24014, -27890, -27838, -31429, -31211, -31087, 
    -31402, -29729, -26847, -23591, -19274, -18566, -13854, -9375, -5826, 
    -2367, 3501, 6362, 11813, 14807, 20375, 21887, 24433, 27136, 30116, 
    29806, 31627, 32208, 30228, 28644, 26873, 25525, 21413, 17678, 14353, 
    11146, 5213, 1959, -2888, -6640, -12023, -13737, -18633, -23153, -24093, 
    -26214, -29803, -30090, -30554, -29822, -29595, -30027, -26943, -24127, 
    -21866, -19638, -16051, -11469, -5931, -1571, 2667, 5968, 11876, 15734, 
    18769, 21602, 24358, 26118, 27566, 31361, 31209, 31367, 30758, 28281, 
    28485, 24556, 22363, 17257, 16219, 10914, 6324, 1165, -3191, -7758, 
    -10695, -14985, -18236, -22721, -23756, -28724, -27708, -30103, -30893, 
    -31746, -31423, -29410, -26742, -22927, -20825, -17920, -15307, -11246, 
    -6060, -2106, 1100, 5082, 11778, 14674, 19668, 20928, 25906, 27129, 
    27089, 29704, 30151, 30295, 29844, 28163, 26418, 24759, 21218, 18065, 
    13368, 10834, 7161, 572, -1073, -7085, -10093, -13242, -17726, -21305, 
    -24339, -27984, -30109, -30231, -30037, -31725, -30224, -28605, -29084, 
    -26069, -22000, -16998, -15887, -11107, -7135, -3050, 1084, 6756, 10130, 
    15196, 18978, 20920, 24263, 27222, 29096, 30520, 31349, 30285, 30182, 
    30186, 27342, 25435, 21199, 18037, 16683, 12175, 6333, 2257, -1886, 
    -6642, -11171, -15101, -17853, -21240, -24703, -26295, -29309, -29636, 
    -30387, -29888, -30778, -29358, -27550, -23415, -22311, -18694, -16950, 
    -11218, -8448, -3314, 1483, 5700, 9108, 15055, 17675, 22649, 23510, 
    26726, 29589, 29907, 30058, 30927, 29788, 28217, 26867, 26469, 22056, 
    19823, 16254, 12776, 7460, 3879, -1187, -4742, -9636, -13973, -18318, 
    -20312, -24542, -26769, -29691, -30356, -32030, -31918, -30548, -28651, 
    -28265, -25340, -23500, -18757, -16356, -12720, -7330, -2667, 2204, 4984, 
    9429, 13442, 17035, 21088, 24317, 27277, 27517, 30109, 29270, 30537, 
    31809, 28212, 27361, 25379, 22578, 18343, 17175, 12329, 8570, 4217, -915, 
    -5749, -9968, -13213, -16004, -19082, -24333, -26803, -27980, -28605, 
    -32206, -30398, -30505, -28962, -27466, -26088, -23072, -18548, -14971, 
    -11689, -9043, -5190, 382, 5068, 8726, 11918, 17242, 21813, 22785, 25451, 
    29716, 29518, 29352, 31959, 30487, 30920, 28053, 25512, 22596, 20908, 
    16532, 13322, 8484, 4343, 1106, -5054, -8818, -12804, -17285, -19012, 
    -23775, -25663, -28943, -29878, -31043, -31329, -30956, -29551, -28421, 
    -25935, -23223, -21711, -17552, -13039, -9935, -5695, -316, 4004, 9152, 
    12892, 17467, 20334, 22447, 27281, 26203, 29670, 30792, 32302, 29722, 
    29649, 28289, 26302, 24538, 20212, 16846, 13690, 8833, 4429, 1785, -5649, 
    -8064, -12073, -15842, -21031, -22709, -24768, -28565, -29576, -31980, 
    -30616, -29737, -29911, -27763, -24666, -24667, -19615, -16652, -13813, 
    -8305, -5827, -302, 4916, 8961, 11824, 17410, 19760, 22422, 25401, 29125, 
    30092, 30622, 29700, 30013, 30877, 28314, 26609, 22800, 19303, 15699, 
    14553, 9774, 5869, 378, -4080, -6941, -12899, -15669, -18786, -24431, 
    -26525, -28785, -29052, -29045, -29902, -30663, -29812, -29499, -25271, 
    -22934, -22030, -17790, -14128, -9905, -5348, -1566, 3562, 7184, 12223, 
    14442, 18860, 22609, 26186, 27646, 28520, 30038, 29587, 30484, 29661, 
    29603, 25652, 23746, 21092, 18206, 13854, 9075, 5177, 1696, -4093, -8301, 
    -11738, -15692, -17639, -23948, -25863, -27450, -28894, -29625, -31509, 
    -31049, -31788, -28415, -26454, -24561, -20235, -16558, -15079, -10621, 
    -5596, -1761, 4571, 7856, 11034, 15849, 19062, 20593, 25911, 27863, 
    28355, 29854, 31042, 32363, 29276, 28863, 27334, 24415, 21268, 17890, 
    15053, 10471, 6799, 1384, -1624, -7837, -11573, -16255, -19158, -22014, 
    -25598, -28224, -28458, -31071, -29982, -29165, -28530, -28946, -25357, 
    -24915, -20597, -18940, -13160, -10731, -7579, -2389, 2200, 8172, 12685, 
    15569, 17369, 21685, 25276, 26161, 30136, 31302, 32092, 30297, 29265, 
    29037, 26600, 25698, 22092, 17902, 13966, 10119, 6325, 1780, -3304, 
    -7123, -11028, -14414, -17776, -20174, -25046, -27611, -27866, -28867, 
    -31334, -30246, -29673, -29558, -26586, -25362, -22254, -19375, -14660, 
    -10216, -6673, -1927, 1431, 7554, 11539, 13225, 18195, 21264, 24022, 
    26776, 28331, 30530, 30635, 30433, 30486, 28450, 28323, 23686, 20456, 
    18698, 14272, 9801, 6221, 2026, -755, -5775, -9516, -13359, -17330, 
    -22158, -24696, -27774, -28538, -29203, -31947, -31581, -28786, -28981, 
    -28420, -23716, -20575, -18176, -15544, -12309, -5312, -3044, 1649, 6521, 
    8870, 15177, 17563, 21614, 24768, 25853, 29022, 30088, 30713, 31029, 
    29982, 28902, 26875, 25768, 22647, 18855, 15313, 10195, 7772, 3257, 
    -1722, -5744, -8986, -12842, -18990, -20192, -23572, -26480, -28380, 
    -28966, -31013, -31438, -31128, -29056, -26975, -24612, -22751, -19985, 
    -14858, -12032, -8652, -2790, 1192, 6994, 9887, 13693, 17839, 21069, 
    24702, 26075, 30188, 28563, 30805, 29841, 30880, 27728, 25983, 25444, 
    23660, 19266, 14968, 11441, 8355, 3567, -1467, -6369, -8374, -13727, 
    -17396, -20683, -24877, -25063, -29108, -29281, -29841, -30679, -31330, 
    -28335, -28647, -25097, -23050, -19143, -15013, -12373, -9072, -2742, 
    1468, 4373, 8637, 12298, 18735, 20166, 24291, 27526, 28700, 29153, 31066, 
    30988, 30452, 28800, 27030, 25244, 22941, 21035, 15927, 13207, 7970, 
    2219, 668, -5780, -8273, -13302, -16747, -21788, -24614, -27112, -28536, 
    -28134, -31677, -30994, -30455, -29786, -26107, -25966, -23283, -20478, 
    -16741, -11830, -8078, -4064, 811, 4352, 9330, 11768, 15535, 19527, 
    23823, 25810, 26833, 30274, 30373, 31914, 29044, 29740, 28524, 26101, 
    24094, 20939, 15914, 12353, 9422, 5298, -225, -4696, -10245, -12725, 
    -16269, -20624, -24022, -26021, -28865, -30993, -30313, -29711, -30209, 
    -29544, -29196, -26109, -22638, -19820, -16447, -11860, -7612, -3044, 
    -450, 4315, 8323, 13097, 16314, 19211, 23376, 25256, 26636, 29274, 30650, 
    31241, 30782, 29997, 28968, 25983, 24398, 20002, 16896, 13672, 8318, 
    3697, 852, -4889, -6912, -13308, -15596, -20970, -23063, -26041, -27992, 
    -28871, -30310, -30666, -29583, -29454, -28284, -27044, -23558, -19943, 
    -17704, -13172, -9605, -4650, -1260, 3355, 8647, 12257, 15896, 21459, 
    22266, 26355, 27702, 29555, 30985, 30293, 30144, 30692, 29242, 25793, 
    23252, 21872, 18210, 12982, 9793, 5006, 826, -4256, -9440, -11341, 
    -16782, -18126, -22172, -24956, -28789, -29329, -30762, -32211, -29767, 
    -30689, -28094, -26276, -24503, -21748, -17904, -14418, -10191, -5423, 
    -1584, 4047, 6844, 11910, 15961, 21303, 23884, 26322, 28335, 29727, 
    29053, 30265, 31112, 30073, 28668, 27016, 24328, 20995, 17025, 14684, 
    9748, 4679, 1083, -2084, -7519, -12835, -15085, -19248, -22535, -24453, 
    -27477, -29702, -30919, -31276, -29813, -29794, -29516, -26713, -24843, 
    -21758, -16828, -13350, -9966, -6043, -738, 4043, 8464, 11299, 15541, 
    19986, 22512, 25008, 28178, 29739, 29809, 30840, 30862, 30151, 30319, 
    26933, 23620, 21392, 18002, 13861, 8657, 7250, 181, -2870, -7533, -9878, 
    -15559, -19452, -21047, -25441, -27773, -27692, -30499, -29846, -30570, 
    -28797, -27479, -27100, -24433, -19821, -17900, -14258, -9163, -6889, 
    -2063, 2680, 6169, 11177, 14605, 18510, 22722, 24482, 26460, 30728, 
    30379, 30262, 30141, 31189, 28325, 26964, 24208, 21923, 19154, 12870, 
    11273, 6237, 1551, -1170, -5158, -9957, -15104, -19257, -21279, -25765, 
    -26357, -28590, -30440, -30277, -29386, -30285, -28714, -28504, -23644, 
    -21449, -18269, -14547, -11105, -7952, -2524, 3263, 7850, 10470, 15239, 
    18400, 21353, 24255, 27545, 28526, 29745, 30759, 31552, 29591, 27767, 
    26907, 25287, 20488, 18621, 14142, 10318, 8282, 1323, -1933, -7040, 
    -9400, -14181, -19126, -21618, -24287, -26029, -27705, -30283, -31083, 
    -30844, -31010, -29223, -25749, -25847, -21238, -18820, -15101, -10583, 
    -7301, -2228, 3174, 5985, 10263, 14547, 18173, 20096, 23782, 26555, 
    30021, 30136, 31820, 29512, 28908, 29065, 28421, 24308, 21635, 18974, 
    16355, 10470, 8193, 2841, -511, -4342, -10069, -13452, -18454, -21401, 
    -25407, -26043, -28269, -29917, -30997, -30772, -29589, -29133, -26505, 
    -26769, -21735, -19114, -15588, -11895, -7813, -2766, 986, 4799, 9479, 
    14571, 18976, 22045, 24479, 25598, 28202, 30199, 30747, 30890, 30932, 
    29404, 28294, 26408, 22301, 19417, 15980, 11088, 8214, 3513, -2013, 
    -5118, -9314, -12862, -16925, -19729, -24660, -26531, -26778, -29867, 
    -31555, -31834, -28845, -30557, -28169, -25704, -23644, -18654, -14147, 
    -12349, -6901, -4101, 1166, 4181, 9832, 14223, 18120, 20000, 23491, 
    26187, 29204, 29311, 30509, 30398, 30175, 29483, 28723, 26144, 22342, 
    19123, 16099, 13682, 7656, 2529, -340, -4947, -9865, -13130, -16396, 
    -20620, -23952, -25618, -27989, -30128, -30479, -30465, -30894, -30117, 
    -28201, -27517, -22349, -20562, -17272, -11558, -8085, -3896, -1160, 
    4501, 8605, 12410, 17643, 21186, 24448, 25072, 28338, 31442, 29625, 
    30244, 31198, 30072, 27676, 25659, 22889, 20124, 17242, 13378, 9539, 
    4216, 1492, -4728, -8816, -13867, -15466, -21157, -23937, -26770, -27339, 
    -29474, -31060, -31481, -30736, -29424, -27236, -25671, -24358, -20223, 
    -17139, -13420, -9749, -5067, -941, 5104, 8446, 12581, 16864, 20986, 
    24424, 25121, 28375, 30990, 30971, 32056, 30473, 30022, 28201, 25178, 
    24267, 19956, 17476, 13191, 7288, 5369, 1622, -3671, -8498, -12142, 
    -18148, -21489, -22740, -25227, -26914, -31102, -30669, -30158, -31728, 
    -28567, -28735, -26580, -23420, -21596, -16072, -13055, -9925, -6386, 
    -1339, 2328, 9185, 13238, 16111, 18918, 23736, 24346, 28220, 29277, 
    30685, 32226, 30780, 29618, 27802, 26589, 23369, 21352, 17816, 14518, 
    9859, 5406, 1374, -2496, -8362, -11293, -15819, -19767, -22923, -26037, 
    -28571, -29301, -29189, -29767, -30457, -29808, -27516, -25824, -23770, 
    -20985, -16498, -13351, -9613, -5164, 670, 2560, 6935, 11502, 14104, 
    18596, 23587, 25819, 28566, 29159, 29909, 30364, 29871, 29565, 28728, 
    26858, 24200, 20029, 17445, 12956, 9957, 4370, 948, -3252, -7110, -12709, 
    -16294, -19247, -23391, -25613, -27532, -27738, -32089, -32379, -31229, 
    -28153, -27889, -25715, -23050, -20449, -19180, -12889, -10764, -4368, 
    -918, 3753, 6321, 12085, 14607, 19416, 21279, 23772, 27352, 29132, 30490, 
    29500, 30026, 29487, 30278, 26460, 24580, 21179, 18167, 13077, 10140, 
    6293, 2417, -3764, -7224, -11976, -15088, -20315, -21502, -24932, -27876, 
    -29039, -30675, -30176, -31906, -29607, -29245, -26087, -24862, -22261, 
    -18039, -13735, -10862, -6583, -1882, 1673, 6943, 10462, 15079, 19440, 
    22443, 24208, 26403, 28648, 30192, 29963, 31553, 29818, 30320, 27663, 
    25696, 22410, 18638, 13563, 11443, 6518, 2515, -2290, -6390, -11087, 
    -15734, -18829, -21492, -25662, -27382, -28770, -29470, -30271, -31608, 
    -29128, -29626, -27269, -24603, -21899, -18772, -14219, -9651, -6527, 
    -2022, 1522, 4917, 10567, 14284, 17764, 21678, 24207, 27858, 29038, 
    29094, 30551, 31673, 29330, 28298, 28381, 25625, 21477, 19807, 15174, 
    11304, 5742, 2429, -739, -6901, -11668, -13692, -16613, -22018, -24885, 
    -26217, -29324, -29362, -31430, -29178, -31793, -29781, -25755, -24941, 
    -22918, -19114, -15772, -12448, -5429, -2421, 1875, 5580, 8961, 13580, 
    16430, 21571, 25718, 26240, 30056, 29667, 31156, 30649, 29950, 27727, 
    27253, 24010, 21574, 18175, 14642, 10653, 6079, 3508, -568, -6097, -8727, 
    -13745, -16889, -21656, -23878, -26353, -29048, -30697, -30443, -29901, 
    -29775, -27983, -27852, -26503, -21211, -20658, -14716, -12592, -6461, 
    -3172, 1403, 4615, 9592, 13830, 15997, 20145, 23616, 27220, 27904, 28579, 
    31015, 31627, 31367, 28500, 28199, 26290, 22555, 19968, 15540, 10844, 
    8593, 4414, -1145, -4803, -8169, -14880, -16298, -21025, -23783, -25686, 
    -27371, -31021, -30896, -31346, -30324, -28946, -28837, -26825, -22776, 
    -19791, -15910, -11285, -6767, -3556, 1293, 5625, 8950, 13796, 16472, 
    21141, 24371, 25113, 28293, 29418, 30371, 30267, 30984, 28419, 27019, 
    26020, 23308, 19825, 17314, 13976, 8389, 3635, -517, -4566, -9854, 
    -13112, -16859, -19541, -23720, -26191, -28512, -31067, -29151, -31062, 
    -31759, -29904, -27575, -25627, -21173, -18546, -15796, -10700, -9411, 
    -4630, 1286, 4168, 7904, 13840, 17749, 20482, 23391, 26519, 27941, 29645, 
    31639, 31093, 31164, 30075, 28587, 25606, 23657, 19842, 15482, 13008, 
    8658, 3438, -550, -3473, -8605, -12592, -17020, -18511, -23252, -25133, 
    -28147, -29576, -29921, -30879, -29101, -28549, -28028, -26679, -24057, 
    -18465, -15064, -13437, -8599, -4536, 1110, 4358, 9489, 13333, 15677, 
    19469, 22725, 24876, 28618, 30380, 30379, 30323, 30436, 29745, 28604, 
    25448, 23831, 20880, 16884, 12472, 8969, 5589, 1030, -4065, -9319, 
    -11921, -16806, -18865, -23405, -26134, -27802, -30280, -29317, -30017, 
    -31859, -29508, -29570, -26549, -23816, -18810, -16294, -12728, -10385, 
    -5965, -548, 3876, 8398, 11467, 17082, 20009, 21054, 25095, 27375, 30165, 
    31021, 31246, 29773, 29135, 27865, 26200, 25384, 21201, 17542, 13747, 
    10579, 4611, 650, -4286, -7570, -12337, -15677, -19373, -24288, -25517, 
    -26390, -29909, -31413, -30368, -29814, -28001, -27531, -25210, -23135, 
    -21111, -18139, -14204, -11086, -4648, -1719, 1813, 7228, 11450, 15411, 
    19328, 22631, 26857, 27687, 29913, 31057, 29964, 30586, 29138, 28583, 
    26666, 23873, 20418, 18882, 13425, 9562, 5842, -246, -4457, -7651, 
    -12786, -14766, -19252, -23187, -24360, -25840, -28079, -30311, -30587, 
    -29264, -28956, -27822, -25493, -24101, -20578, -17825, -13503, -9233, 
    -5569, -1069, 2170, 6947, 10628, 16460, 19778, 22416, 24933, 26763, 
    29560, 29957, 31754, 30333, 28929, 28265, 25079, 24349, 21035, 18220, 
    12867, 8938, 6084, 1606, -3060, -6075, -11290, -15708, -17356, -20942, 
    -25518, -25563, -27952, -29629, -30378, -31455, -31617, -28985, -27166, 
    -25587, -21344, -17986, -15111, -10238, -4668, -2331, 3210, 6617, 11497, 
    14990, 18708, 21826, 24570, 25707, 30094, 29877, 29996, 29243, 30428, 
    28654, 25750, 25284, 21724, 18181, 15595, 8889, 6778, 1785, -2741, -6700, 
    -10713, -14112, -17690, -22942, -25282, -27106, -29590, -31362, -31407, 
    -30913, -30211, -28088, -27353, -23043, -21071, -18455, -14813, -10154, 
    -6006, -1702, 1942, 6497, 10832, 15579, 17278, 20673, 23352, 25588, 
    27320, 30001, 29338, 30785, 30594, 28641, 27713, 25328, 21765, 18164, 
    14503, 10127, 7303, 3419, -3187, -5223, -11391, -14936, -17914, -21213, 
    -23013, -27648, -29638, -31077, -30899, -29837, -28683, -29019, -27256, 
    -24339, -21323, -18250, -15652, -11033, -6389, -2985, 1946, 4843, 11688, 
    14120, 17147, 22209, 23649, 26908, 28451, 30164, 31434, 31887, 30731, 
    28348, 28455, 25689, 21127, 18898, 13559, 12868, 5516, 2835, -322, -7199, 
    -10094, -15265, -19714, -21663, -23510, -25618, -27337, -29124, -31280, 
    -31576, -28716, -27961, -27705, -25273, -22885, -18047, -15209, -11490, 
    -7682, -2041, 1311, 3935, 9606, 13794, 18588, 20218, 23231, 26640, 29348, 
    28113, 31861, 30187, 31712, 28838, 27144, 24256, 23949, 20714, 15957, 
    11448, 7558, 3819, -1533, -3795, -11107, -12866, -18275, -21293, -24290, 
    -26831, -27094, -30696, -28927, -30715, -29902, -30436, -27144, -26382, 
    -21545, -21209, -16707, -11378, -8237, -4843, -481, 3966, 9471, 13377, 
    16210, 20591, 24817, 26441, 28196, 29924, 30154, 30785, 30644, 29404, 
    29323, 24795, 22087, 19349, 15712, 11764, 8004, 4231, -582, -6333, -8682, 
    -13285, -17525, -20873, -22806, -25810, -27983, -28853, -30619, -30859, 
    -30393, -29984, -27865, -26904, -21867, -19724, -17280, -13025, -8385, 
    -5166, -65, 6141, 8814, 12542, 17479, 21587, 23760, 26778, 28991, 30751, 
    29647, 31139, 30675, 30188, 27792, 26196, 22888, 20735, 15942, 13261, 
    8406, 5417, 376, -5522, -8811, -14084, -16680, -20625, -22196, -26505, 
    -27298, -28871, -29637, -29853, -31926, -28121, -27198, -27023, -24244, 
    -21474, -16148, -11342, -8678, -5514, 185, 5591, 7845, 12763, 16082, 
    18912, 22454, 26397, 27028, 28152, 30981, 30736, 30849, 30431, 27714, 
    26825, 24009, 20297, 15590, 13728, 10074, 5616, -636, -5033, -8758, 
    -12923, -16734, -20254, -23927, -24572, -28504, -28372, -30970, -30771, 
    -29787, -29525, -26649, -26694, -24092, -19662, -17465, -13540, -10538, 
    -3578, -499, 5188, 7359, 11953, 17274, 19990, 22880, 27134, 28909, 29084, 
    29023, 30559, 31061, 30150, 28460, 26398, 22710, 20646, 17025, 13643, 
    8331, 4528, 738, -5011, -8142, -12211, -17718, -19493, -22855, -27128, 
    -28280, -29010, -30341, -30044, -30471, -29934, -27950, -26894, -23191, 
    -19097, -18085, -14622, -9617, -4409, -2164, 3570, 6120, 12170, 16070, 
    20840, 22557, 24641, 27348, 31158, 30684, 32070, 30655, 29332, 30245, 
    27407, 22742, 19621, 17621, 14172, 9582, 5446, 1407, -3594, -8880, 
    -10654, -16423, -19102, -22210, -24348, -27373, -29247, -30640, -31363, 
    -30955, -29809, -27636, -27504, -24020, -20207, -17215, -12281, -11028, 
    -5904, -1631, 4112, 7513, 13267, 15802, 19402, 23595, 25829, 27968, 
    28650, 31417, 31820, 30460, 30585, 28629, 26326, 23250, 21185, 18334, 
    14702, 11000, 7210, 1846, -2785, -7801, -12763, -16304, -18507, -21862, 
    -23787, -28346, -29256, -29722, -30897, -31497, -29014, -27657, -27575, 
    -24584, -22972, -18766, -14443, -10079, -6136, -194, 1980, 6246, 9936, 
    15067, 18639, 21855, 25012, 28973, 29723, 32069, 29181, 30423, 29612, 
    27940, 27655, 24668, 20556, 18182, 15703, 10787, 5356, 1072, -1203, 
    -5332, -11667, -14505, -19719, -22620, -24894, -26018, -30474, -30033, 
    -30224, -29489, -29797, -28985, -28054, -25376, -21621, -18635, -16253, 
    -10418, -5330, -2091, 1837, 5682, 11561, 15584, 19451, 20855, 24281, 
    25594, 30379, 29957, 31640, 30672, 30462, 28968, 28321, 24434, 21897, 
    17983, 15287, 10207, 8367, 846, -2880, -6880, -11258, -14680, -18146, 
    -21289, -23209, -27552, -27868, -29308, -30296, -31284, -30504, -29597, 
    -27221, -25180, -21201, -17762, -14449, -11562, -6412, -1790, 2003, 7463, 
    9162, 14002, 16990, 21899, 24208, 25721, 28746, 30859, 30464, 30116, 
    29220, 29766, 26878, 23860, 22481, 19682, 14995, 11225, 8705, 1623, 
    -1269, -5249, -9961, -14998, -19168, -21782, -24727, -26390, -27980, 
    -29234, -29787, -29526, -31464, -28770, -28248, -25120, -23530, -20094, 
    -16395, -12468, -8245, -2861, 1446, 6487, 9820, 14613, 17848, 21470, 
    23815, 26160, 29163, 29400, 32231, 30425, 30227, 29859, 28308, 26754, 
    23570, 19399, 15368, 11730, 7787, 3838, -676, -6338, -10250, -14149, 
    -18251, -21424, -25785, -27196, -26597, -31014, -31693, -31495, -29682, 
    -29916, -27849, -25427, -23361, -19413, -14621, -11708, -9077, -4301, 
    475, 4837, 10419, 14367, 17925, 21767, 23925, 27293, 28287, 29785, 29635, 
    29777, 30740, 30075, 28915, 25892, 21394, 19393, 14943, 13864, 7451, 
    2885, -1232, -4750, -9227, -13940, -16552, -21093, -22583, -24646, 
    -27765, -29453, -30999, -29643, -31531, -28375, -28694, -26573, -22509, 
    -21583, -16260, -13935, -8522, -4835, 934, 3828, 7781, 14607, 16695, 
    19346, 22255, 25864, 27926, 29114, 32051, 31687, 30351, 28004, 27941, 
    25924, 22882, 20135, 16513, 12444, 8681, 3037, 80, -4624, -9105, -12656, 
    -15608, -20278, -23132, -25458, -28268, -28908, -30014, -30910, -30918, 
    -28813, -29027, -25074, -25044, -20689, -16618, -13544, -10047, -3788, 
    87, 5307, 8352, 12883, 15478, 20510, 23579, 26708, 27944, 29353, 29538, 
    30017, 30220, 30468, 28988, 26943, 24007, 21591, 17370, 12036, 7919, 
    5618, 155, -4003, -8759, -12515, -16419, -20409, -22762, -26215, -27896, 
    -30603, -28957, -30166, -30715, -30087, -28282, -25314, -23241, -20333, 
    -15980, -13791, -10320, -4451, -452, 2740, 8233, 11780, 15202, 21219, 
    22184, 24868, 28402, 29401, 30199, 30438, 29868, 30514, 29267, 26978, 
    22604, 22084, 16544, 12461, 8449, 4466, 1381, -3015, -9353, -12064, 
    -15114, -20891, -22880, -24694, -28512, -30093, -30607, -30786, -31630, 
    -30036, -29329, -26586, -24845, -20428, -17463, -13337, -8493, -4244, 
    145, 4841, 7705, 11698, 15618, 19559, 22726, 24112, 27335, 30271, 30983, 
    30567, 29318, 30568, 29763, 27904, 24900, 22502, 17679, 13246, 9889, 
    6170, 1380, -2840, -8802, -10724, -14665, -19510, -21042, -23931, -27768, 
    -28873, -29910, -30727, -31281, -28806, -27578, -26190, -24438, -20054, 
    -17599, -14699, -10132, -4872, 178, 2387, 7794, 12877, 14058, 17999, 
    23658, 25854, 27737, 30048, 28824, 30755, 28809, 30127, 29368, 25313, 
    24320, 20295, 17809, 13686, 10834, 5124, 1720, -3189, -6428, -9913, 
    -15694, -17221, -22920, -25099, -26946, -28947, -31267, -30468, -29581, 
    -30703, -27789, -26874, -25841, -20776, -18766, -13703, -10252, -7383, 
    -2934, 2525, 8270, 11100, 15339, 19342, 21556, 25321, 26593, 28112, 
    29331, 30745, 31902, 30444, 28216, 27062, 24521, 20493, 17018, 14395, 
    10981, 4737, 2520, -2237, -8117, -10798, -15552, -19537, -21681, -24753, 
    -27590, -27898, -29395, -31721, -30736, -29077, -28336, -27290, -26125, 
    -22675, -16833, -14738, -9892, -7714, -3714, 2382, 7121, 10395, 13979, 
    18294, 20802, 24779, 26735, 28850, 29742, 29757, 30627, 29018, 28634, 
    26613, 25019, 20956, 19876, 14455, 10855, 5125, 2401, -2858, -6676, 
    -10568, -15646, -18942, -20634, -24239, -26693, -29977, -29527, -30796, 
    -30164, -30517, -29255, -26536, -25370, -22826, -18473, -15355, -11779, 
    -6341, -1536, 1048, 5366, 10002, 14819, 17819, 21373, 24824, 26837, 
    29342, 30538, 29960, 30932, 31094, 27785, 26440, 23814, 22406, 18853, 
    15871, 11024, 5853, 1852, -1864, -7392, -10870, -13718, -16702, -21376, 
    -24022, -27920, -28554, -31186, -31886, -31065, -30986, -29137, -27224, 
    -25266, -23960, -20057, -14703, -10660, -6736, -4324, 1334, 5548, 8327, 
    12303, 17796, 21729, 24977, 26472, 27941, 29081, 31692, 31025, 29569, 
    29298, 27902, 25357, 22440, 20035, 15865, 10841, 8198, 4147, -1102, 
    -5484, -11159, -14089, -17907, -20185, -24339, -26110, -29827, -29933, 
    -29737, -32313, -29334, -30281, -27413, -24278, -22244, -20098, -14668, 
    -11327, -8502, -3568, 1366, 3924, 10317, 14017, 16797, 21193, 23742, 
    24844, 28482, 30254, 30131, 30318, 31059, 29131, 28390, 26665, 22647, 
    19752, 16197, 12537, 7209, 4123, -1550, -4855, -8390, -13131, -15383, 
    -20455, -22458, -27229, -28477, -29314, -29751, -30456, -29669, -28775, 
    -28527, -26942, -22755, -18561, -15666, -12138, -6794, -2320, -735, 5472, 
    9057, 13187, 15318, 19890, 24033, 26830, 28448, 29422, 30927, 30100, 
    30964, 30097, 27740, 26255, 21631, 21545, 16422, 11203, 8551, 5636, 162, 
    -4290, -8842, -14375, -16812, -20363, -22068, -26084, -28463, -29970, 
    -29667, -31896, -30577, -28386, -28242, -26411, -24331, -20565, -14862, 
    -12351, -7806, -4772, -702, 3442, 9669, 13158, 16587, 20181, 24502, 
    25183, 28036, 29864, 30347, 29866, 30777, 30639, 28293, 24836, 23117, 
    21533, 16410, 11511, 9860, 5471, -807, -3578, -9342, -11059, -15995, 
    -20431, -21791, -25300, -27408, -28965, -30928, -30599, -30396, -29671, 
    -27454, -26372, -24374, -19164, -18496, -14124, -9735, -4426, 51, 3121, 
    8000, 10612, 17168, 19798, 23989, 26985, 27080, 30584, 31877, 30893, 
    29675, 30631, 28665, 25499, 24114, 20525, 16414, 14797, 8857, 5934, 555, 
    -4274, -8105, -11934, -17062, -19941, -23607, -25659, -26735, -29289, 
    -31056, -30961, -31023, -29306, -28023, -26498, -24100, -19456, -15794, 
    -13307, -9522, -3786, -396, 4288, 7707, 11278, 14552, 20074, 23539, 
    27105, 27309, 29192, 29291, 31593, 31136, 30832, 28668, 25662, 23980, 
    22025, 16662, 13427, 8994, 5580, 1680, -3201, -8328, -13126, -14490, 
    -19642, -22331, -24683, -28651, -28501, -30140, -30373, -30566, -29601, 
    -27100, -27862, -22640, -20401, -17537, -14090, -10045, -5437, -1713, 
    4581, 7700, 10240, 14306, 18103, 22110, 23950, 28292, 28156, 30049, 
    30141, 31615, 29928, 27947, 26001, 23292, 20040, 18405, 13824, 9088, 
    6929, 1739, -1966, -6673, -11291, -14388, -19126, -22790, -25432, -27837, 
    -27269, -30037, -31407, -31985, -31002, -29449, -27133, -25226, -20457, 
    -17352, -12992, -10340, -5530, -1007, 2355, 6594, 12527, 15299, 17894, 
    21503, 25015, 26787, 28941, 29619, 30491, 32017, 28865, 29925, 27265, 
    24148, 21388, 18643, 14321, 9960, 8171, 2687, -1407, -7531, -11451, 
    -15488, -18581, -22490, -24389, -26913, -28691, -30159, -31178, -30902, 
    -30939, -29145, -26831, -24647, -21754, -19567, -16407, -9894, -7172, 
    -2708, 1019, 6663, 10474, 13933, 17668, 21093, 24721, 27259, 29526, 
    30023, 30443, 31237, 28851, 27804, 26563, 24189, 22813, 19933, 15559, 
    10870, 7974, 2048, -2384, -6674, -10015, -13916, -19069, -21990, -25128, 
    -27118, -28371, -29589, -30615, -31047, -28968, -28693, -26633, -25956, 
    -23098, -18984, -13936, -11480, -7134, -1731, 1214, 7606, 9184, 13682, 
    18095, 21793, 24532, 26666, 27280, 28728, 30567, 30830, 30838, 28918, 
    26819, 25651, 20655, 20242, 16804, 11275, 5928, 2712, -1192, -6485, 
    -11367, -14293, -19427, -22161, -25226, -25332, -28332, -29669, -30631, 
    -29133, -30450, -29474, -26808, -25016, -21228, -19978, -14369, -10885, 
    -6323, -2095, 2215, 5653, 8759, 14717, 18344, 19821, 23440, 27874, 27172, 
    30392, 31016, 31462, 30600, 30045, 28202, 26453, 23935, 19842, 15646, 
    12147, 6382, 2812, -1043, -6399, -9912, -14118, -17506, -19971, -23116, 
    -27116, -28046, -31265, -30688, -31295, -31310, -30458, -28276, -26398, 
    -22278, -19198, -16107, -12377, -7165, -3015, 932, 3841, 9339, 12774, 
    17504, 21341, 23509, 27359, 28118, 28954, 31715, 30781, 30851, 29137, 
    28815, 26353, 22222, 17970, 15012, 12866, 8199, 4533, -676, -5502, -9569, 
    -13894, -17773, -20316, -23481, -27197, -27662, -30548, -31787, -31153, 
    -30459, -29348, -27295, -24844, -22632, -19793, -14974, -13565, -7577, 
    -2951, 111, 4312, 9857, 13087, 17451, 21649, 23262, 25725, 28289, 30071, 
    32073, 30553, 31470, 30740, 26844, 24828, 23018, 20697, 16064, 11559, 
    7628, 4965, -973, -5622, -8751, -14128, -17974, -21126, -23691, -25435, 
    -27793, -28885, -30172, -31115, -31055, -28082, -28153, -26087, -23309, 
    -20916, -16407, -12135, -9026, -4137, 518, 5968, 8228, 12705, 15517, 
    20803, 22262, 26075, 27969, 30290, 32156, 29689, 28977, 29547, 28039, 
    26263, 22549, 21061, 18408, 12688, 8449, 3955, 1555, -3227, -9156, 
    -12833, -15751, -20333, -22104, -25762, -27868, -29610, -31001, -29176, 
    -30595, -29110, -27165, -25391, -23438, -21279, -17055, -13054, -9528, 
    -4024, -1539, 3576, 8834, 11521, 16103, 19318, 23238, 24137, 28065, 
    30733, 31420, 30389, 31060, 30410, 27442, 27141, 24674, 21507, 17845, 
    12803, 10285, 5634, -564, -3194, -7557, -13223, -15726, -19439, -22985, 
    -25914, -28847, -29429, -29423, -31486, -28974, -30229, -28278, -27394, 
    -23959, -21269, -15974, -12942, -8803, -4651, -1619, 3858, 8155, 11125, 
    14595, 19218, 22095, 25091, 26166, 28920, 30859, 32144, 29808, 28954, 
    27567, 26087, 24314, 20846, 17280, 14961, 9999, 5866, 1122, -1982, -7504, 
    -12474, -15707, -17855, -22441, -25120, -28652, -29782, -31044, -30398, 
    -29257, -29606, -28053, -27585, -24012, -21651, -18579, -14103, -10013, 
    -5066, -311, 4221, 7095, 11235, 15794, 18767, 22676, 24942, 25729, 29520, 
    28827, 31096, 28874, 30630, 28886, 25635, 25398, 22093, 17671, 13476, 
    10400, 6405, 3040, -2366, -8191, -12311, -16688, -19377, -22092, -24526, 
    -27801, -29219, -30103, -29658, -31166, -29338, -28341, -27264, -25613, 
    -20825, -17735, -13739, -10340, -5849, -3278, 2035, 7317, 11482, 14910, 
    18379, 21905, 26395, 27291, 29377, 29978, 30543, 31275, 30369, 29525, 
    27701, 25247, 22350, 18227, 15139, 10967, 7210, 1915, -3407, -5484, 
    -10702, -13902, -19734, -21810, -24186, -27752, -29896, -30899, -29285, 
    -30888, -29794, -30008, -27660, -23239, -22283, -18092, -15067, -11469, 
    -6363, -2362, 1523, 7041, 10741, 15009, 18253, 21644, 25073, 26963, 
    27297, 30406, 29613, 32568, 28693, 28396, 26601, 25725, 21628, 18075, 
    15250, 9750, 6031, 2748, -2554, -7016, -11476, -13641, -17913, -20746, 
    -24456, -27790, -28991, -28877, -32270, -31072, -30271, -27156, -26438, 
    -25017, -23105, -18163, -15569, -11137, -6387, -3807, 2671, 4177, 9898, 
    14832, 17492, 20618, 24417, 28050, 29473, 29499, 30856, 30971, 29848, 
    29745, 26875, 26373, 21453, 19358, 13968, 12541, 7215, 2986, -2133, 
    -5038, -11149, -13610, -18289, -22724, -23974, -26285, -28100, -31098, 
    -32379, -29951, -30124, -29033, -28322, -25806, -22401, -20073, -15186, 
    -12656, -6284, -2543, 1286, 6717, 10210, 13592, 16596, 21438, 24828, 
    26906, 29150, 29659, 29888, 31242, 29739, 27823, 27554, 24865, 23013, 
    18215, 16619, 12441, 8690, 3399, -768, -4143, -9513, -12945, -17651, 
    -20725, -23946, -26335, -27576, -28577, -31544, -30371, -30396, -29950, 
    -27035, -25457, -22437, -20389, -15262, -11590, -9584, -3627, 258, 5724, 
    9260, 13368, 17549, 21551, 23988, 25536, 28566, 29681, 29783, 32461, 
    30577, 27965, 29299, 24728, 22855, 20512, 16052, 11667, 7851, 2937, -838, 
    -4804, -9101, -12982, -18022, -20751, -23229, -26319, -27188, -29368, 
    -30584, -29875, -30103, -30225, -26606, -26184, -22489, -20836, -16048, 
    -12079, -8589, -5272, 891, 4199, 10019, 13232, 17564, 21205, 22520, 
    26189, 29310, 29343, 29750, 30907, 31715, 30266, 27417, 25093, 21705, 
    20183, 17243, 11797, 6990, 2811, -867, -4879, -9258, -12685, -16611, 
    -21467, -23581, -26521, -29188, -29948, -32014, -30714, -30765, -28448, 
    -28178, -26544, -22903, -20105, -16613, -12555, -9310, -3751, -427, 4635, 
    8046, 12583, 17920, 19295, 23344, 25492, 28032, 29584, 28840, 32166, 
    29745, 28326, 27745, 25515, 23088, 21784, 16720, 13222, 10450, 6210, -66, 
    -3528, -8510, -12337, -17643, -19579, -23770, -26493, -28294, -29842, 
    -29788, -30902, -31714, -29791, -27002, -25613, -23795, -21656, -15272, 
    -13317, -10267, -4621, -487, 3894, 9294, 12111, 16742, 20344, 22747, 
    25581, 27195, 28344, 31128, 31640, 31671, 30822, 27032, 26402, 23688, 
    19783, 16498, 14153, 9649, 3920, 539, -3703, -7391, -11884, -15523, 
    -19606, -21920, -24859, -27389, -29224, -30595, -31308, -29790, -29530, 
    -29385, -25691, -24253, -20646, -18233, -12923, -8958, -5280, -1331, 
    3089, 6633, 10311, 16850, 19647, 22385, 25300, 27877, 29504, 30966, 
    31512, 30704, 30125, 29779, 27038, 24592, 20149, 18067, 14929, 10351, 
    4158, 348, -3441, -7895, -11722, -15411, -18860, -22233, -25427, -26519, 
    -28982, -30934, -31564, -31147, -30107, -29287, -25804, -23960, -20500, 
    -17676, -12877, -8838, -7152, -1420, 3437, 8334, 11237, 15635, 19012, 
    23263, 26485, 27894, 29956, 30803, 31958, 30145, 28740, 27678, 26981, 
    24580, 22555, 17862, 14093, 8953, 5564, 981, -3201, -5612, -11986, 
    -15405, -18181, -22781, -24383, -25979, -29289, -29699, -30361, -30543, 
    -29495, -28158, -27324, -23359, -20816, -18882, -14968, -11222, -5049, 
    -916, 1580, 5851, 10359, 13878, 18703, 21214, 24188, 27223, 29526, 29345, 
    31581, 31789, 28317, 29069, 27010, 24551, 21576, 17778, 13689, 10999, 6622, 
    3676, -2026, -5695, -12381, -14487, -19561, -23188, -23177, -27932, 
    -28690, -29536, -32057, -29969, -31467, -30009, -28441, -24307, -21274, 
    -17311, -15270, -9627, -6164, -1596, 1938, 7162, 11031, 14369, 18602, 
    21295, 25589, 27103, 28738, 30627, 31257, 31644, 29856, 29629, 27594, 
    25678, 20945, 19669, 16301, 10389, 6840, 2317, -1944, -6263, -10508, 
    -15123, -18396, -23103, -24469, -26859, -29486, -29000, -30431, -30547, 
    -31050, -29193, -26866, -23443, -22194, -18947, -16075, -11795, -6790, 
    -1442, 1357, 7463, 9393, 14214, 16958, 20624, 23713, 26725, 28047, 29269, 
    29716, 30684, 31476, 29210, 26934, 25089, 24053, 19331, 15775, 10814, 
    7426, 3195, -1232, -5610, -10429, -14669, -17646, -21156, -24630, -25765, 
    -28058, -28798, -31831, -30765, -29642, -29756, -26928, -25470, -23597, 
    -18345, -15015, -11684, -6466, -3298, 479, 4056, 9869, 14130, 16401, 
    19865, 23128, 25225, 28511, 30228, 30293, 29586, 29580, 28750, 28179, 
    24710, 21996, 19483, 16616, 11753, 7601, 3453, -1740, -6019, -8361, 
    -12845, -17170, -22166, -24230, -25649, -27067, -28799, -32112, -31005, 
    -29225, -30305, -27723, -23885, -22822, -18002, -16035, -12478, -7045, 
    -2657, 1023, 4933, 9086, 13677, 17842, 20642, 24364, 25186, 28112, 29191, 
    29717, 30747, 31201, 30602, 28704, 25983, 21945, 18879, 15953, 13402, 
    8193, 4049, -1164, -4452, -9983, -13838, -17194, -19570, -23480, -25190, 
    -26754, -29413, -31043, -30806, -29009, -30733, -27276, -24960, -22342, 
    -19035, -15599, -11186, -8363, -5079, 641, 3820, 10403, 11812, 17735, 
    20504, 23367, 25897, 27287, 29430, 29719, 30102, 28933, 28639, 28326, 
    26055, 22570, 20421, 16130, 11410, 8933, 4715, 593, -3169, -9340, -13348, 
    -18332, -21107, -23963, -24804, -28378, -29568, -29657, -30481, -30331, 
    -29712, -29161, -25555, -22530, -20148, -16567, -12921, -8290, -5204, 
    897, 5290, 8815, 12789, 16549, 21018, 24101, 25861, 28165, 28983, 28728, 
    29833, 31740, 28989, 27312, 25151, 23964, 19331, 15435, 12497, 9115, 
    6239, 398, -5271, -7113, -11386, -16310, -20560, -23109, -27290, -26495, 
    -29074, -32013, -31290, -30395, -28506, -28191, -26403, -22672, -20949, 
    -17333, -12598, -9089, -5167, -813, 2720, 8385, 12164, 17020, 19839, 
    23427, 24824, 27468, 28756, 30574, 31154, 31144, 29457, 27782, 25668, 
    23446, 19977, 17768, 14612, 9762, 4448, 2064, -2967, -7987, -11962, 
    -16571, -18560, -22731, -25371, -28924, -29505, -29928, -32201, -30082, 
    -29433, -27738, -26448, -24412, -19933, -18882, -14034, -10665, -4294, 
    -368, 2415, 8111, 11425, 16074, 19761, 22729, 25289, 26433, 28474, 31323, 
    30496, 31054, 29556, 28821, 26911, 24521, 21140, 18502, 13816, 11373, 
    5119, 731, -3250, -6857, -11591, -14412, -18641, -22513, -24682, -28607, 
    -29764, -30965, -31030, -30600, -28999, -28346, -27387, -24025, -20718, 
    -16853, -14599, -10113, -6810, -1779, 2564, 6751, 10792, 15739, 19808, 
    23486, 23868, 28573, 27963, 30889, 30774, 30479, 30351, 28855, 25173, 
    23958, 22160, 17078, 12606, 9277, 5333, 1783, -1587, -6598, -11597, 
    -16399, -19864, -21762, -24532, -26499, -29884, -30536, -29950, -30611, 
    -30922, -28504, -27028, -24613, -23236, -17356, -13604, -9552, -4764, 
    -1445, 2773, 7135, 11240, 14087, 19452, 22382, 25432, 27243, 29896, 
    30561, 30755, 31006, 29911, 27542, 26921, 25578, 20828, 19375, 14172, 
    11800, 7414, 2343, -2730, -7185, -11486, -13692, -17723, -21632, -24354, 
    -27715, -29499, -29201, -29838, -29679, -30526, -27860, -26751, -25453, 
    -21209, -20255, -15417, -10813, -6124, -2052, 1481, 6406, 12130, 15157, 
    18425, 21444, 23762, 27706, 28463, 30048, 29520, 30208, 29948, 29142, 
    26525, 24440, 20500, 18250, 14207, 11311, 5151, 3365, -3148, -5010, 
    -10573, -14162, -17169, -22018, -22922, -26525, -28734, -29067, -30912, 
    -30261, -30687, -28951, -27793, -23505, -23465, -20440, -15524, -10635, 
    -7006, -3633, 649, 7155, 10331, 15076, 18027, 22183, 24455, 25948, 28630, 
    29851, 30417, 30087, 30303, 27885, 26262, 25477, 23137, 18248, 15564, 
    11139, 6462, 1820, -1161, -6287, -10086, -14736, -17012, -20868, -23857, 
    -26799, -29603, -30673, -31943, -30461, -31073, -27793, -26052, -25125, 
    -23251, -19275, -16242, -11880, -7157, -2871, 240, 6685, 10490, 14863, 
    18033, 21165, 24593, 27829, 27995, 29284, 30944, 31450, 28781, 29791, 
    26661, 24763, 21847, 19061, 15203, 13152, 6993, 3769, 228, -4018, -9931, 
    -15051, -18080, -21764, -24124, -26023, -28137, -28426, -31863, -30874, 
    -31468, -30188, -26850, -25205, -22448, -19070, -15714, -11924, -8410, 
    -2633, 1950, 5220, 9555, 13358, 17024, 20666, 23030, 26922, 27313, 29827, 
    31556, 31666, 30214, 29306, 28047, 25251, 22091, 19833, 15946, 10642, 
    7936, 3909, -283, -5974, -9841, -12153, -18307, -20601, -24424, -25056, 
    -28413, -29834, -29949, -30279, -31698, -29671, -29059, -25693, -23230, 
    -19957, -16830, -12895, -7809, -4479, -1165, 5863, 8041, 13249, 16088, 
    21322, 24345, 24640, 28870, 28276, 30417, 31688, 29773, 30146, 27696, 
    24818, 23542, 19131, 18269, 11874, 10024, 5444, -266, -4873, -9044, 
    -13182, -17981, -21915, -24474, -26726, -27895, -28585, -30349, -31480, 
    -30096, -28691, -27211, -25426, -22169, -21161, -15232, -11038, -8709, 
    -3598, -569, 4346, 9120, 12992, 16241, 20158, 22888, 26537, 28541, 28842, 
    31232, 30880, 30784, 30674, 28180, 25227, 22840, 20240, 15538, 12559, 
    8984, 4506, 185, -5368, -8384, -13537, -15792, -20704, -22710, -27121, 
    -28543, -30594, -29621, -32156, -30221, -29171, -27690, -26018, -22296, 
    -20796, -16987, -11827, -9044, -5635, -1067, 5513, 7527, 11892, 17287, 
    19758, 23268, 26485, 26800, 29508, 29234, 31115, 30953, 30179, 27711, 
    25010, 23615, 20418, 15945, 14532, 9968, 5154, -476, -4920, -7078, 
    -10541, -15075, -19722, -22280, -24878, -27009, -29982, -30023, -31688, 
    -30597, -29411, -28510, -26540, -22345, -21982, -17847, -14444, -9499, 
    -5095, -1563, 2359, 7127, 12705, 16174, 19486, 21473, 25322, 29528, 
    29272, 29737, 32600, 31423, 28818, 29455, 25521, 22728, 21068, 19259, 
    12833, 8411, 6708, 1109, -2342, -7754, -11749, -14982, -18111, -21968, 
    -25101, -28652, -28330, -31898, -30718, -30450, -29226, -28705, -28454, 
    -23953, -21960, -18007, -14282, -10533, -5080, -1502, 3223, 8850, 12143, 
    16573, 19802, 22432, 25708, 28886, 29063, 31194, 31150, 29820, 29039, 
    28986, 26735, 23214, 19910, 16421, 15330, 11261, 6124, 1652, -2938, 
    -6401, -10679, -13810, -17998, -23185, -26298, -27060, -29134, -30449, 
    -31208, -32068, -29749, -28490, -27371, -23824, -21138, -17888, -13648, 
    -11806, -6398, -2045, 2077, 5901, 12228, 14599, 18345, 22134, 24553, 
    28425, 28304, 31102, 30544, 30276, 30672, 28431, 28446, 23432, 20172, 
    17785, 15221, 11051, 7672, 2452, -2771, -6147, -11662, -14753, -19934, 
    -21850, -23340, -26813, -28851, -30471, -31126, -30036, -29837, -27980, 
    -26717, -25788, -22873, -20254, -13574, -10164, -4934, -1846, 2797, 5694, 
    9800, 15173, 19099, 20313, 24387, 26876, 28747, 29494, 31053, 31614, 
    29419, 28797, 27036, 23211, 21795, 16782, 15537, 11981, 6859, 2667, 
    -2543, -6255, -10429, -14657, -18804, -22180, -24511, -25909, -27888, 
    -30498, -31305, -30112, -30727, -30267, -26601, -24211, -22111, -17259, 
    -13851, -11712, -7003, -3059, 2094, 6622, 10819, 14847, 17795, 21025, 
    24807, 26741, 28118, 29963, 31094, 30566, 28488, 29527, 27355, 25624, 
    21871, 19119, 14263, 10782, 6893, 3776, -2546, -7140, -10221, -12682, 
    -19663, -21791, -24346, -27831, -28460, -30730, -31113, -31652, -31471, 
    -29443, -26764, -24816, -21710, -18787, -15506, -11326, -6316, -4203, 
    1142, 7358, 9174, 13299, 17871, 21056, 23167, 26820, 26869, 30532, 32293, 
    32304, 30268, 27647, 26871, 26621, 22381, 21010, 16207, 12113, 7472, 
    3812, -1979, -6169, -11110, -13633, -17132, -20608, -23592, -24969, 
    -29041, -29809, -30431, -31913, -30674, -28254, -26162, -27102, -23981, 
    -19110, -15986, -11533, -8080, -3258, 1150, 4008, 9715, 12679, 18793, 
    21180, 22548, 25950, 26674, 31482, 30445, 31332, 29494, 28010, 28503, 
    25557, 21880, 19929, 15211, 12357, 8621, 4734, -693, -5598, -9584, 
    -12333, -16104, -20546, -24405, -27187, -27089, -29842, -30208, -30836, 
    -30678, -30984, -26876, -26715, -22709, -20360, -16501, -12712, -8873, 
    -3173, 409, 4287, 8048, 12586, 17449, 21365, 23689, 26226, 28443, 31075, 
    31260, 30737, 31168, 29782, 27702, 25494, 24201, 19067, 16709, 12089, 
    8220, 3747, -1415, -5459, -10244, -13473, -15977, -19850, -22123, -26789, 
    -28075, -30246, -29564, -30478, -30560, -29047, -28828, -26048, -22891, 
    -19587, -16225, -13501, -8110, -4252, 558, 4267, 8708, 14266, 16854, 
    19403, 24226, 26033, 27901, 28522, 28700, 31833, 31091, 29920, 28200, 
    27226, 23347, 21581, 17022, 12493, 8752, 3597, 1111, -2746, -8842, 
    -11118, -16792, -19575, -22815, -26115, -27797, -27928, -31201, -31060, 
    -29333, -29810, -28839, -25910, -24004, -21562, -16732, -13656, -10279, 
    -4819, 709, 3524, 7865, 12683, 16883, 18752, 23245, 26205, 28176, 30397, 
    29467, 31070, 30869, 30046, 28106, 26660, 22880, 20449, 17167, 13274, 
    9987, 4858, -517, -4703, -8851, -11481, -16112, -18896, -22427, -24851, 
    -26280, -29583, -31723, -31367, -31583, -29563, -27981, -25448, -23220, 
    -20952, -17158, -13453, -10161, -4286, -1142, 4226, 6644, 11407, 16145, 
    18413, 23438, 25958, 28583, 29326, 30363, 30069, 29128, 29237, 28856, 
    27299, 23731, 20916, 16734, 13932, 8911, 5530, 978, -3730, -7424, -11462, 
    -16113, -20622, -21405, -25277, -26587, -29520, -31880, -29648, -30264, 
    -29715, -29670, -26452, -24921, -21935, -17675, -15597, -9647, -4792, 
    -1355, 1995, 6453, 11749, 15365, 19802, 21089, 26132, 26515, 28836, 
    30154, 29637, 31671, 29929, 28130, 26947, 23181, 19662, 17002, 14571, 
    8941, 5970, 115, -1350, -7089, -10715, -15622, -19691, -22314, -24445, 
    -26383, -28783, -31766, -30824, -30789, -30159, -28532, -26464, -23499, 
    -21365, -17578, -13937, -9754, -7474, -1869, 3462, 7737, 11162, 14408, 
    19549, 22791, 24164, 26629, 28865, 31213, 31045, 31989, 29740, 27803, 
    25321, 25013, 20439, 17727, 14278, 9166, 5569, 3106, -1587, -6569, 
    -12553, -16216, -19390, -22106, -24280, -25499, -29473, -30370, -30874, 
    -30924, -30894, -28922, -27942, -25498, -21552, -19701, -15762, -10923, 
    -7288, -2469, 2539, 6277, 10819, 14665, 19279, 22816, 26073, 28171, 
    28262, 29046, 31007, 30184, 30277, 27853, 27279, 23934, 21988, 19297, 
    14838, 12577, 6718, 1351, -2856, -7632, -11714, -15244, -16927, -22366, 
    -24715, -26229, -29581, -29512, -30839, -30298, -30257, -28926, -28470, 
    -23684, -22190, -19784, -14020, -11852, -7760, -3273, 2849, 4563, 9147, 
    13180, 19383, 20788, 24896, 27366, 28751, 30451, 29771, 29983, 29946, 
    29443, 28085, 26404, 21038, 18542, 14257, 10460, 6616, 2724, -2029, 
    -6874, -9848, -14845, -18673, -22566, -25074, -26318, -28018, -30484, 
    -31893, -30695, -31393, -28189, -26982, -24044, -22456, -19628, -14453, 
    -10745, -7060, -3795, 790, 5202, 10400, 13778, 18106, 21409, 25325, 
    27075, 28689, 30405, 30958, 31425, 31776, 27856, 27326, 26305, 22586, 
    19630, 15329, 12977, 8040, 2141, -916, -5485, -10078, -12041, -18941, 
    -21561, -23989, -26068, -28166, -29246, -30888, -30993, -31744, -28435, 
    -26624, -24693, -21669, -19374, -16571, -12900, -7882, -2497, 1163, 5755, 
    9433, 12441, 16019, 20078, 25061, 26561, 28007, 29250, 31179, 30804, 
    31373, 28230, 28747, 24822, 22477, 19200, 16256, 11207, 8246, 4089, 
    -1570, -3943, -10140, -12633, -16195, -19570, -23700, -28128, -28345, 
    -29576, -30010, -30385, -30504, -28671, -28343, -26377, -24307, -19966, 
    -16499, -11556, -8381, -4640, -732, 4772, 9022, 13303, 16075, 19111, 
    22910, 26292, 26818, 30001, 30575, 29863, 29608, 29722, 27934, 26497, 
    22539, 20159, 16289, 12580, 8768, 3891, -143, -3039, -7636, -12533, 
    -18071, -20670, -23181, -26130, -28287, -29525, -31340, -32041, -30721, 
    -28618, -26939, -25951, -24154, -20297, -16119, -13934, -9147, -5281, 
    -554, 3446, 7555, 11100, 15426, 20181, 22505, 26437, 27442, 29284, 31175, 
    30882, 31248, 30557, 26734, 25107, 23865, 19743, 17038, 13611, 9158, 
    5386, -656, -5377, -9691, -12633, -15793, -20195, -21458, -24891, -28335, 
    -29714, -29986, -31758, -30239, -28764, -28949, -27848, -21940, -20646, 
    -17179, -11405, -8996, -5879, 91, 4844, 7605, 13981, 16212, 20130, 21934, 
    24892, 28168, 29216, 30907, 31292, 31426, 30675, 29671, 25959, 25431, 
    20395, 17433, 14929, 10004, 5105, -89, -3756, -8081, -12770, -15440, 
    -19847, -21427, -26136, -27179, -28521, -29073, -30387, -30608, -30889, 
    -28295, -26868, -24073, -20779, -15856, -14267, -9021, -6048, -445, 4860, 
    6536, 13314, 14426, 19913, 24265, 24500, 28189, 29337, 30724, 31401, 
    30769, 29959, 28242, 24961, 24159, 20730, 17940, 14428, 9580, 5085, 732, 
    -3083, -7354, -12031, -15270, -19968, -22479, -24394, -27853, -29418, 
    -29935, -31210, -30940, -29378, -27089, -26454, -24321, -20485, -17269, 
    -15120, -9362, -5566, -2316, 2143, 8001, 11354, 15565, 17513, 22314, 
    24283, 26209, 29712, 31509, 29982, 30635, 29911, 29417, 27992, 24244, 
    19626, 18444, 13524, 9776, 5785, 1368, -1960, -6763, -11452, -14642, 
    -20064, -21413, -24806, -28671, -29357, -28658, -31957, -30008, -30199, 
    -29732, -26342, -24888, -22538, -19368, -14891, -10348, -4903, -3135, 
    1689, 7671, 11474, 16719, 17861, 21797, 23748, 28308, 29679, 30516, 
    31020, 31705, 28981, 29227, 27079, 24582, 21761, 17596, 15178, 11775, 
    6282, 1585, -1951, -7972, -11400, -13684, -17901, -23525, -24439, -28255, 
    -29011, -28618, -30940, -30803, -29589, -29719, -28193, -24906, -20589, 
    -18681, -14387, -10221, -6229, -3238, 2404, 5712, 11798, 15389, 18919, 
    21251, 24801, 28086, 29993, 30920, 30555, 30199, 31021, 28637, 28502, 
    25169, 21295, 17509, 15594, 11299, 5935, 2653, -1800, -5746, -11379, 
    -13474, -18750, -21144, -23277, -27158, -27971, -28271, -29763, -29994, 
    -30110, -28024, -28112, -24989, -22535, -18505, -16042, -11153, -7154, 
    -1738, 1683, 5158, 10025, 13943, 18714, 22547, 25379, 27154, 28649, 
    31444, 30241, 31048, 29947, 29491, 26049, 23285, 21979, 18239, 14854, 
    10800, 7485, 2319, -1857, -6340, -10317, -14740, -17973, -21271, -24021, 
    -26082, -30128, -30786, -30700, -29281, -30025, -28650, -29074, -26419, 
    -21910, -18138, -16420, -12106, -6601, -2739, 1426, 5914, 9687, 13862, 
    17931, 21497, 24255, 25973, 27875, 31051, 30978, 29521, 30815, 29970, 
    26217, 24753, 21820, 17631, 15414, 11793, 8027, 2895, -1201, -5558, 
    -9269, -13172, -17077, -21195, -22657, -26542, -28172, -30855, -30654, 
    -29727, -30624, -28842, -28595, -24995, -24148, -18149, -14778, -11929, 
    -7278, -4594, 1930, 4100, 10398, 13374, 18195, 21294, 23443, 25871, 
    28992, 31204, 29954, 31215, 29623, 29284, 28259, 25546, 22493, 18424, 
    14291, 12480, 6980, 3318, -1084, -4222, -8818, -12710, -16974, -21540, 
    -22841, -26164, -29398, -29197, -31185, -30471, -30440, -29210, -28241, 
    -24817, -22837, -20299, -16259, -10975, -8922, -3223, 1104, 4518, 9257, 
    12411, 17875, 20182, 24241, 26702, 28722, 29879, 30809, 30758, 31475, 
    29941, 27047, 24006, 22747, 19351, 16134, 12698, 9690, 4333, 840, -4696, 
    -8851, -12100, -17532, -20364, -23549, -26152, -29500, -28100, -31490, 
    -29866, -29668, -30737, -28088, -25317, -23078, -20184, -18095, -13205, 
    -7864, -5629, -945, 5425, 9550, 13137, 15205, 20063, 22833, 25929, 28615, 
    30614, 31923, 30827, 31350, 27847, 27123, 24820, 22973, 21281, 18602, 
    12527, 7208, 5406, 283, -4018, -8867, -13323, -15677, -21331, -22763, 
    -25607, -27684, -29411, -31618, -30986, -31176, -30332, -27492, -26303, 
    -24526, -19781, -17671, -13264, -10671, -5068, 202, 4198, 7594, 12295, 
    16753, 19013, 22856, 26984, 26498, 29721, 29764, 29597, 29366, 31112, 
    27098, 24993, 25398, 21226, 16683, 14317, 10034, 5042, 851, -3036, -8733, 
    -11080, -15650, -21014, -23608, -26087, -28670, -29105, -30326, -32083, 
    -30361, -28526, -28307, -25678, -24354, -21065, -17177, -15066, -9416, 
    -5243, -586, 2499, 8227, 12413, 16209, 20851, 24204, 25718, 28838, 30208, 
    29547, 31014, 31938, 29731, 28836, 26558, 24086, 19460, 16273, 14503, 
    9418, 4514, 866, -2462, -8023, -11899, -16409, -19984, -21500, -24949, 
    -27647, -29851, -31193, -31120, -30727, -29889, -28841, -27398, -24587, 
    -22042, -17109, -14033, -9907, -6147, -1294, 3216, 8738, 13161, 15508, 
    18925, 22955, 23612, 27589, 29945, 30123, 31274, 31090, 30907, 28681, 
    27428, 25533, 22264, 18075, 14369, 10136, 7193, 1104, -3278, -7743, 
    -10982, -15089, -18857, -20966, -24772, -26870, -28788, -31748, -30798, 
    -30824, -30309, -28042, -26569, -24366, -21050, -19945, -14715, -9862, 
    -5934, -1782, 2979, 7562, 9973, 16259, 18316, 22528, 24928, 27133, 28787, 
    29744, 30070, 29913, 29725, 29531, 27298, 24093, 20873, 18537, 14774, 
    10262, 7710, 2323, -1795, -6746, -12298, -14801, -18700, -21842, -23791, 
    -25482, -29105, -30542, -30469, -31087, -30049, -28209, -26125, -24373, 
    -21535, -18779, -13973, -10622, -7156, -3601, 1737, 6669, 9643, 14615, 
    18635, 22926, 25616, 26003, 29385, 29451, 31640, 30628, 29869, 29159, 
    27227, 25493, 20458, 18068, 14294, 9640, 7811, 2299, -759, -6386, -10277, 
    -13528, -19977, -21498, -24327, -25395, -28793, -30851, -30183, -31460, 
    -31711, -30427, -28756, -23963, -21774, -19476, -15711, -11847, -7936, 
    -2498, 149, 5677, 10511, 13118, 17773, 23129, 23097, 25354, 27779, 30090, 
    31725, 29906, 28898, 29374, 26817, 25168, 23923, 17089, 14641, 12010, 
    8420, 2094, -1497, -5955, -8944, -14836, -18111, -21456, -24209, -27935, 
    -29318, -29298, -29404, -31437, -29004, -28537, -27337, -24606, -22579, 
    -18605, -15019, -10589, -7249, -2792, 385, 7166, 9322, 14581, 19003, 
    21050, 23638, 27200, 26843, 30813, 31248, 31227, 30206, 29192, 26704, 
    24972, 22998, 19419, 15869, 13069, 7044, 4072, -2388, -4419, -10397, 
    -13846, -17003, -20857, -24230, -25145, -29221, -30235, -30079, -30590, 
    -30945, -28856, -28918, -26047, -21870, -18791, -15821, -10580, -6783, 
    -3100, 620, 3991, 9571, 13550, 16245, 20778, 23965, 26360, 27852, 30980, 
    30072, 29519, 29261, 31100, 26690, 26100, 23817, 19561, 15008, 13297, 
    6347, 3595, 247, -6546, -9660, -12820, -17793, -22113, -22482, -26545, 
    -27937, -29506, -30514, -31539, -30209, -27639, -28641, -24895, -23343, 
    -19289, -15990, -12541, -7452, -3903, 704, 4984, 9912, 14471, 17701, 
    19892, 23473, 25237, 27400, 29632, 29995, 30315, 30440, 29345, 27282, 
    25380, 23433, 20663, 15843, 12821, 8647, 5482, -901, -6186, -9403, 
    -11978, -17795, -21469, -22783, -26148, -28143, -29804, -29395, -29784, 
    -30267, -29824, -26929, -25353, -22318, -20642, -16249, -12788, -8369, 
    -3944, -450, 3826, 9582, 12446, 16537, 19628, 24320, 26712, 29387, 30288, 
    29487, 31482, 30346, 28843, 28801, 26672, 24710, 20850, 16857, 13528, 
    9905, 3090, 1204, -3078, -7974, -12454, -15782, -21439, -22214, -26309, 
    -28883, -29299, -30357, -29308, -30235, -29391, -29630, -25185, -25073, 
    -20108, -17929, -12017, -10153, -4903, -161, 3767, 7505, 12398, 17452, 
    18996, 23222, 26586, 27350, 29738, 29577, 31672, 29786, 30566, 28045, 
    26460, 23529, 20476, 16153, 12979, 8804, 3528, 2296, -2653, -7340, 
    -11970, -15788, -18457, -22458, -25134, -28896, -30174, -29502, -31443, 
    -29669, -29105, -29258, -25463, -24013, -19251, -17274, -12910, -9031, 
    -6812, -1389, 3009, 6738, 12732, 14138, 20087, 24186, 24935, 29088, 
    27718, 31517, 30529, 31654, 28066, 30029, 26217, 22704, 21103, 17856, 
    13330, 9487, 5744, 1422, -2716, -7900, -10726, -15861, -18243, -22191, 
    -25764, -26527, -30186, -30631, -30056, -29940, -29615, -27498, -27228, 
    -23820, -20321, -17783, -12430, -8912, -5922, -1232, 2927, 6778, 11851, 
    14882, 19268, 23499, 25352, 26358, 28309, 30057, 30342, 30579, 30791, 
    28152, 26755, 24046, 20108, 18579, 14250, 10222, 7276, 1527, -2006, 
    -7692, -11904, -14787, -20522, -23576, -24755, -27925, -28287, -29866, 
    -30539, -30273, -28775, -27113, -26659, -25343, -21216, -17740, -13987, 
    -10614, -4716, -1294, 4123, 7037, 12254, 15180, 19306, 23430, 23953, 
    26294, 29210, 31481, 29435, 31190, 30480, 28547, 26016, 23824, 22307, 
    18673, 15062, 11001, 6652, 3693, -1435, -5957, -11048, -15414, -17874, 
    -21725, -24275, -28502, -28801, -29910, -30435, -30102, -31164, -28228, 
    -26310, -23581, -22560, -17649, -14867, -11304, -6832, -1062, 2020, 5943, 
    10507, 14583, 17631, 22086, 25138, 25980, 29949, 30379, 30630, 30985, 
    31260, 27338, 27989, 25222, 21926, 17452, 14446, 10955, 7219, 2842, 
    -1967, -7183, -11161, -12919, -18361, -19940, -25339, -27914, -28595, 
    -31457, -29669, -29960, -28940, -28982, -25428, -25577, -21686, -18486, 
    -15506, -12202, -6685, -3416, 3334, 5385, 10098, 13614, 17496, 22244, 
    23797, 27345, 29901, 28660, 31727, 29837, 30651, 28198, 25928, 25066, 
    22957, 19571, 15511, 11084, 6895, 4333, -1007, -6229, -9151, -12710, 
    -18129, -20161, -23492, -26098, -28064, -28995, -29635, -30925, -29822, 
    -28610, -26319, -24126, -22634, -18436, -15649, -13150, -6743, -3120, 
    1239, 6921, 10441, 14075, 19161, 22190, 23979, 26293, 27749, 30781, 
    29092, 31321, 29227, 28335, 27788, 25309, 22120, 19575, 16747, 10716, 
    8817, 3147, -960, -4999, -9958, -13823, -17233, -21667, -24395, -27574, 
    -28973, -30413, -30800, -30652, -29197, -29062, -27590, -24392, -23323, 
    -19896, -14876, -11582, -8116, -3038, 599, 5516, 10962, 15011, 16470, 
    19689, 24030, 26643, 30185, 30685, 30505, 31833, 32042, 29263, 28747, 
    24607, 22414, 18956, 16115, 11195, 6230, 3394, -762, -4345, -10096, 
    -14197, -18481, -20282, -22981, -26787, -28933, -28483, -30823, -29617, 
    -31307, -29350, -27598, -24422, -22646, -19398, -15572, -11653, -9367, 
    -5557, -58, 4202, 8884, 13991, 18156, 19337, 22612, 26354, 27089, 29396, 
    30562, 30647, 30106, 29584, 27916, 24952, 22864, 19445, 16584, 13312, 
    7714, 4298, 422, -4251, -8855, -14487, -17023, -21659, -23902, -26988, 
    -27994, -29229, -30900, -30064, -30095, -30086, -28381, -25261, -22208, 
    -19476, -16644, -12530, -9732, -4470, 154, 4929, 8146, 13736, 18182, 
    20012, 24250, 24631, 28403, 30694, 30316, 29730, 29995, 28951, 29026, 
    26168, 23344, 19682, 15649, 12264, 9425, 5133, -974, -4467, -8359, 
    -12636, -15709, -20060, -23610, -24603, -27969, -30221, -30959, -31560, 
    -29416, -28779, -26462, -26024, -22733, -21524, -17473, -14615, -8913, 
    -4617, -905, 4743, 8445, 12741, 16095, 19329, 23005, 24696, 28630, 28574, 
    31150, 31152, 30467, 29611, 27015, 25732, 25009, 21122, 17663, 13523, 
    9655, 5793, -86, -3720, -8263, -12548, -15651, -20393, -22051, -25192, 
    -28345, -28505, -29219, -30923, -30698, -29242, -29439, -27211, -22896, 
    -21098, -16473, -14611, -9315, -5011, -675, 3155, 7362, 10914, 17452, 
    19531, 22606, 26319, 27182, 29189, 30133, 32065, 29716, 29660, 29120, 
    25907, 24424, 19842, 16559, 13243, 11183, 4910, 1510, -3266, -6769, 
    -11875, -15069, -19922, -23201, -26852, -28515, -29048, -30007, -30398, 
    -30795, -30108, -28311, -26756, -24466, -21221, -17969, -12752, -10988, 
    -5823, -2146, 3196, 7861, 12827, 16306, 19313, 23021, 25650, 28819, 
    29535, 30399, 30848, 30182, 29454, 28842, 26760, 24694, 21209, 16922, 
    15086, 11545, 5281, 1833, -3190, -7963, -11639, -14419, -19595, -22481, 
    -23554, -26612, -28377, -30691, -30780, -30049, -31287, -28628, -26261, 
    -24339, -22825, -18134, -14639, -10943, -6124, -1260, 2238, 5845, 11029, 
    16034, 18765, 20192, 24295, 28069, 28708, 29691, 30823, 31212, 31677, 
    28002, 26496, 24724, 20999, 17675, 13538, 12187, 5204, 2088, -3039, 
    -8256, -10825, -14267, -18398, -21856, -24485, -26598, -27864, -30466, 
    -30857, -31132, -31248, -29651, -28005, -24537, -21506, -18640, -14188, 
    -10729, -5984, -2037, 1821, 6385, 11616, 14728, 19918, 20791, 26220, 
    26172, 28958, 29803, 29895, 29023, 31208, 29169, 27109, 25497, 21018, 
    18598, 15613, 11646, 6806, 2012, -1032, -4680, -9221, -15571, -17874, 
    -20176, -25314, -28352, -30003, -29911, -29277, -30573, -30567, -29244, 
    -26615, -25216, -22281, -19427, -15891, -10894, -7133, -3006, 1385, 4492, 
    8816, 13404, 17116, 21529, 24472, 26198, 28467, 29957, 31069, 31714, 
    29786, 29531, 27905, 24189, 20922, 18572, 15420, 11802, 6402, 4440, 
    -1505, -7587, -10739, -14630, -19397, -21474, -24639, -26004, -27412, 
    -29099, -30787, -32177, -30155, -29280, -28405, -25925, -21774, -19705, 
    -14819, -9809, -6319, -3562, 1273, 6201, 9588, 14010, 17970, 21019, 
    24337, 27627, 29205, 29437, 31100, 29098, 30734, 29855, 28247, 25302, 
    23154, 19187, 16821, 12009, 7692, 1897, -1481, -5199, -9731, -12105, 
    -16057, -22375, -23422, -26217, -27284, -30067, -31571, -29810, -29970, 
    -29832, -28494, -25406, -21984, -19468, -15981, -12713, -8607, -3046, 
    -596, 4471, 11117, 15011, 19162, 19491, 25191, 26328, 26797, 29734, 
    30056, 30061, 29311, 29323, 27877, 24110, 21835, 20069, 16759, 12451, 
    7262, 3523, -1034, -4488, -8903, -12842, -18118, -21380, -22962, -26113, 
    -27752, -30059, -32318, -29570, -30155, -29732, -29170, -25765, -23171, 
    -19534, -17253, -12067, -8090, -4204, -877, 5144, 8891, 12321, 16698, 
    19944, 23247, 27620, 27125, 30364, 30658, 29493, 29806, 29629, 26740, 
    24570, 22288, 19574, 17226, 11185, 8749, 3199, -552, -4492, -8529, 
    -14482, -16719, -20857, -23374, -24745, -27769, -30802, -30340, -31592, 
    -28777, -29516, -27679, -25485, -23038, -20139, -16086, -13119, -7998, 
    -5423, 1017, 3810, 8214, 13332, 17663, 19129, 23543, 27767, 27452, 30038, 
    31314, 29119, 31029, 30793, 28239, 27635, 23127, 18869, 17329, 12341, 
    9310, 3549, 1541, -3159, -9803, -12130, -16123, -19788, -24478, -27265, 
    -27762, -28848, -29728, -31812, -31705, -29034, -27796, -26505, -22259, 
    -21947, -16735, -13299, -10163, -5195, 77, 3019, 7988, 11620, 16489, 
    21347, 22269, 26080, 28156, 29290, 30319, 30662, 30768, 28458, 28353, 
    26820, 23138, 21643, 16519, 14429, 8930, 4489, 840, -4684, -6965, -13218, 
    -15904, -20627, -23296, -24323, -28835, -29681, -30570, -30014, -29952, 
    -29457, -28597, -26255, -24635, -21725, -16566, -13186, -10815, -5038, 
    -2088, 3723, 9302, 11673, 17369, 20658, 21681, 24871, 28443, 28742, 
    31531, 30444, 29740, 30097, 29577, 26635, 23786, 21669, 17344, 13691, 
    9530, 4870, 1842, -4007, -7158, -12048, -15000, -19140, -23689, -26369, 
    -28549, -29329, -30333, -30619, -29954, -29915, -29220, -25718, -24144, 
    -22109, -18136, -12439, -10471, -5194, -1046, 4027, 7975, 12316, 15397, 
    19558, 23111, 25026, 27377, 28790, 30098, 31011, 31192, 29971, 27149, 
    27459, 25402, 20980, 17997, 14748, 9696, 5587, 1271, -2890, -6059, 
    -11446, -14316, -19984, -21231, -24581, -26930, -29456, -31573, -32268, 
    -29938, -30444, -30259, -26311, -25522, -22419, -18425, -13959, -10698, 
    -6609, -1627, 3258, 6050, 11056, 14123, 17994, 21475, 25008, 28350, 
    28853, 30764, 30874, 30278, 30204, 27819, 27456, 22885, 22301, 19908, 
    15481, 10583, 4449, 1995, -1222, -6747, -11889, -13959, -17838, -23523, 
    -24198, -27122, -29635, -30670, -29584, -29804, -31567, -27852, -27269, 
    -24496, -21610, -19933, -14955, -11361, -5632, -1316, 1694, 5302, 9854, 
    13495, 19384, 22586, 25164, 27475, 29988, 30696, 29331, 30183, 30293, 
    29299, 27862, 24246, 22916, 17392, 14771, 11623, 8024, 1203, -460, -6023, 
    -10812, -14882, -19754, -22429, -25857, -26800, -27882, -28451, -28997, 
    -31774, -30437, -29643, -27379, -25454, -21729, -18946, -14031, -12256, 
    -6696, -1370, 1724, 6115, 10709, 14782, 18686, 21120, 25742, 26804, 
    29263, 30972, 28848, 32467, 31685, 28328, 28089, 25897, 21675, 17874, 
    13907, 9624, 8031, 3357, -1731, -4545, -10191, -13209, -19494, -21222, 
    -22965, -27577, -27508, -31569, -30095, -29880, -31093, -28467, -27223, 
    -24602, -22128, -19546, -16820, -11326, -6330, -2828, 756, 5845, 8814, 
    13370, 17145, 22809, 24422, 25639, 29181, 30107, 29181, 30829, 30188, 
    30247, 28098, 24394, 23567, 20843, 15570, 12941, 5831, 3500, -2481, 
    -5771, -9055, -14492, -16975, -21367, -24824, -27396, -28891, -29099, 
    -30750, -31009, -31871, -30935, -28003, -26653, -21936, -18966, -14893, 
    -11150, -6815, -3061, 1132, 6432, 10484, 14383, 17181, 19492, 23070, 
    24985, 29136, 30676, 30731, 31592, 29301, 28897, 26426, 25743, 22422, 
    19609, 16494, 12393, 7283, 5071, 565, -5683, -10090, -13483, -18828, 
    -19544, -23885, -27004, -29539, -29886, -30840, -29820, -30795, -30160, 
    -28913, -25069, -23019, -20625, -15685, -12303, -8921, -2486, 131, 5973, 
    9790, 14781, 16719, 21980, 24283, 25697, 29977, 29929, 31586, 30944, 
    29712, 28806, 29348, 25066, 21996, 20111, 15202, 11960, 7391, 4184, 
    -1752, -4374, -9237, -11293, -16074, -20689, -23720, -25275, -28491, 
    -30389, -30558, -32701, -31450, -29487, -26951, -25553, -21772, -20455, 
    -16549, -13038, -9066, -3995, 844, 3414, 7465, 12180, 16699, 20539, 
    23585, 26096, 28382, 29330, 29904, 30556, 29985, 29958, 28514, 26603, 
    23549, 20321, 17298, 12327, 9448, 4532, 1946, -4513, -9105, -13617, 
    -16732, -18485, -22804, -26658, -27349, -29685, -31216, -31722, -31858, 
    -29772, -28850, -25322, -24706, -20909, -16223, -13348, -8568, -5130, 
    -741, 2750, 7935, 11250, 16413, 18738, 24427, 25000, 28227, 30021, 31642, 
    31351, 30644, 29573, 28566, 26295, 22626, 22236, 16968, 13393, 10663, 
    4583, 2265, -4465, -7592, -11964, -16711, -21027, -22083, -25791, -27890, 
    -29366, -30660, -29559, -31320, -30774, -28552, -25907, -23716, -20203, 
    -18989, -13657, -9820, -6238, -3, 3147, 8109, 12124, 16115, 20153, 23578, 
    26135, 28152, 29749, 30588, 30648, 29996, 29228, 27678, 24973, 22869, 
    21987, 16843, 12414, 8669, 5666, 1026, -3561, -8382, -11993, -15890, 
    -18691, -23322, -25649, -26271, -28144, -30843, -31899, -29980, -29143, 
    -27888, -27010, -24309, -19513, -17980, -14040, -10981, -5558, -1449, 
    2180, 7045, 11931, 17236, 18490, 21274, 24630, 28072, 28995, 30667, 
    30520, 31142, 29825, 28677, 25525, 24069, 20851, 18246, 15237, 9502, 
    5987, 2009, -3973, -6649, -11815, -15251, -18544, -22106, -25086, -27181, 
    -30509, -30356, -32546, -30811, -30474, -28614, -26657, -23783, -20981, 
    -17798, -13882, -8943, -6423, -2010, 2457, 7362, 11686, 16257, 18313, 
    21182, 24094, 27433, 28883, 30829, 30075, 30974, 29976, 28311, 27626, 
    23328, 20222, 18708, 14037, 9809, 5793, 3120, -1392, -6366, -9946, 
    -16427, -19017, -20759, -24334, -27354, -28676, -29070, -30100, -30431, 
    -30774, -28809, -27693, -24878, -22269, -18780, -14002, -10551, -7471, 
    -2021, 2222, 6449, 11003, 15599, 18346, 20138, 24054, 26867, 28574, 
    28901, 30892, 30116, 29714, 29355, 27813, 25460, 21940, 18737, 15080, 
    9689, 8192, 3649, -1483, -5028, -9829, -13988, -18072, -20370, -25180, 
    -26802, -27773, -31358, -31530, -31783, -29516, -29480, -27258, -24647, 
    -21352, -19232, -15355, -11264, -6937, -3075, 1035, 6624, 10131, 12642, 
    17636, 20748, 24404, 25476, 29960, 28818, 30289, 30680, 29845, 28886, 
    26848, 25702, 22274, 18359, 13546, 11428, 7791, 3240, -1826, -4158, 
    -11278, -13454, -17999, -21094, -23840, -24952, -26829, -30330, -30968, 
    -32027, -31491, -28051, -28125, -25190, -23742, -20073, -16290, -11241, 
    -7439, -4420, 2982, 7315, 9527, 13526, 17317, 20156, 23544, 25397, 28265, 
    29895, 31598, 31603, 30811, 29440, 26883, 24971, 22950, 19023, 14486, 
    11925, 6095, 4278, -1560, -6670, -8191, -12881, -17070, -20965, -25705, 
    -27041, -29364, -29518, -31724, -32307, -29729, -27880, -29153, -25438, 
    -22955, -18348, -16112, -12476, -7650, -3742, 4, 6470, 8982, 13437, 
    18028, 19728, 23797, 26174, 29368, 29207, 30643, 29335, 31059, 30199, 
    28129, 25203, 22226, 21122, 16379, 12113, 8902, 4075, 147, -5018, -10118, 
    -14086, -17244, -21056, -23638, -25661, -29250, -30039, -29956, -30512, 
    -31672, -28831, -27882, -25089, -22316, -20609, -15255, -12504, -8033, 
    -4261, 1361, 5373, 10108, 13310, 16814, 20617, 24677, 26410, 27776, 
    29324, 30874, 31640, 30764, 29383, 26989, 24204, 22989, 19094, 15587, 
    12316, 7677, 4044, -674, -4804, -7907, -12963, -16799, -19451, -23410, 
    -25616, -28100, -29903, -29875, -32006, -31391, -28054, -27506, -27079, 
    -22241, -19899, -17871, -12253, -7380, -4789, 440, 3246, 8643, 12745, 
    17171, 20820, 23464, 24935, 28801, 29991, 30813, 32042, 29236, 30034, 
    29261, 27512, 22873, 19348, 16141, 12907, 9013, 4810, -586, -4171, -7912, 
    -11691, -17061, -19298, -22979, -26457, -27923, -29666, -30328, -29754, 
    -28949, -29005, -26826, -26949, -23567, -19843, -17433, -12667, -9538, 
    -3944, -658, 4997, 7656, 12155, 17228, 19490, 23038, 25386, 27503, 29074, 
    30440, 30425, 29610, 29769, 27853, 26726, 23315, 20790, 17678, 12581, 
    9216, 4695, 1629, -4786, -8319, -13905, -16010, -17931, -23342, -26908, 
    -28127, -28809, -29327, -31579, -30814, -29603, -28205, -25987, -25538, 
    -22298, -17777, -13780, -9232, -6719, -14, 3166, 6920, 10521, 16843, 
    20793, 21766, 24727, 27967, 28820, 31282, 31778, 31385, 29476, 28614, 
    27889, 24540, 20113, 16484, 13892, 11124, 5511, 2610, -1915, -7120, 
    -12610, -15975, -19790, -22380, -23931, -26897, -28474, -31015, -29592, 
    -29371, -28341, -28494, -27412, -24251, -21338, -17734, -14289, -11437, 
    -4387, -1399, 2204, 7371, 12399, 14546, 17808, 22311, 24635, 27085, 
    28032, 30159, 30842, 30267, 29875, 29036, 26897, 23929, 20505, 17719, 
    14707, 9383, 6188, 1286, -2221, -6623, -11593, -16280, -18725, -20869, 
    -23965, -26953, -28824, -31756, -30364, -31515, -30893, -27948, -25228, 
    -25243, -21020, -19561, -13529, -10399, -5394, -847, 3347, 7295, 11115, 
    15617, 18743, 20545, 24889, 27032, 29321, 29954, 31258, 31110, 29517, 
    27551, 25257, 23629, 22370, 17992, 14705, 10182, 7595, 1392, -3146, 
    -6839, -10412, -14129, -17733, -21177, -23516, -28189, -28858, -30010, 
    -31170, -31369, -29992, -27964, -28570, -25409, -20622, -20344, -15901, 
    -9971, -6487, -2845, 2630, 5794, 10328, 14434, 18200, 21162, 24058, 
    27812, 28371, 28518, 31188, 29294, 30094, 28483, 25899, 24069, 21339, 
    18573, 15596, 9729, 7156, 1826, -1942, -7096, -9296, -13769, -18056, 
    -22576, -23307, -28565, -28628, -28929, -29741, -30124, -30508, -27360, 
    -26274, -24602, -21721, -19472, -16336, -11389, -7105, -4002, 2027, 5797, 
    10154, 15193, 18529, 19785, 23577, 27086, 27977, 30399, 29824, 30478, 
    29586, 30925, 26582, 24766, 21337, 18650, 14988, 11061, 6557, 2069, 
    -1315, -6206, -10659, -12798, -18512, -20928, -25402, -27426, -28087, 
    -29721, -30636, -29166, -30286, -28855, -25798, -26048, -22182, -20734, 
    -15402, -11252, -6741, -2415, 638, 4886, 10264, 15227, 17614, 21500, 
    23578, 25355, 28290, 30894, 31482, 30992, 30477, 28838, 28342, 26580, 
    21915, 19794, 15335, 11275, 7353, 3231, 6, -5065, -9413, -14256, -17226, 
    -22452, -24992, -25443, -28335, -29397, -30702, -29507, -30652, -28551, 
    -28496, -23623, -22261, -19378, -15468, -11656, -6701, -3693, 986, 5103, 
    10577, 15041, 17597, 20042, 24063, 26758, 28219, 30687, 29753, 30792, 
    29990, 28116, 27920, 25731, 22575, 20181, 16848, 13487, 7990, 4726, 
    -1271, -5847, -9062, -13899, -17768, -21048, -24047, -26945, -27545, 
    -28704, -32250, -29773, -29894, -29227, -28671, -24620, -23444, -18789, 
    -17347, -11356, -8433, -4113, 1177, 4757, 7564, 14257, 17518, 19245, 
    23630, 27738, 28314, 28652, 30063, 32327, 29276, 30156, 29134, 24790, 
    24655, 20039, 15739, 11126, 8140, 4351, -668, -3914, -9099, -13248, 
    -18248, -20830, -24071, -27231, -29011, -28886, -29481, -30495, -30839, 
    -30770, -28706, -24409, -23874, -20460, -17419, -12998, -8484, -3407, 
    -1730, 5301, 7571, 12900, 17176, 20979, 23573, 26580, 27304, 29693, 
    30914, 31130, 30449, 30460, 28504, 27672, 23042, 20737, 15604, 12539, 
    8647, 5640, 657, -5465, -8469, -13679, -16470, -20252, -23234, -25600, 
    -28336, -28953, -30412, -31128, -29472, -30837, -29368, -26284, -23990, 
    -20264, -16918, -13314, -9471, -4462, 847, 4136, 8542, 12215, 16596, 
    20358, 23697, 26664, 27896, 28788, 29912, 31210, 31202, 30391, 29533, 
    26329, 22639, 21459, 16931, 12655, 9070, 5326, 1476, -4876, -9488, 
    -11013, -15572, -20043, -21767, -25280, -28292, -29229, -30672, -29474, 
    -31280, -29885, -28419, -26800, -24863, -20777, -16141, -13247, -10171, 
    -5693, -1625, 4375, 6548, 13027, 16944, 17971, 21545, 25590, 28462, 
    29538, 31258, 30778, 30585, 30910, 29299, 25868, 25192, 21233, 17777, 
    14672, 8582, 5546, 1622, -3329, -8669, -11949, -16529, -19978, -21994, 
    -26053, -26945, -29592, -30554, -31334, -29165, -30850, -29394, -26889, 
    -23145, -22691, -16926, -14974, -9688, -5602, -1923, 2808, 7630, 11699, 
    15148, 19952, 22801, 25225, 27852, 29161, 29416, 30849, 30424, 29763, 
    27894, 28335, 25373, 20454, 17858, 14347, 10328, 6149, 749, -2662, -7447, 
    -12122, -15051, -18073, -23049, -25175, -27681, -28168, -31185, -31482, 
    -30472, -29590, -29502, -27880, -23989, -22557, -17837, -15496, -10185, 
    -5848, -859, 2580, 8088, 11134, 15507, 20084, 22049, 25700, 27785, 30241, 
    29243, 29707, 30406, 29792, 27639, 25760, 23839, 21937, 18251, 14889, 
    9693, 6232, 2423, -1647, -5909, -9645, -14494, -18045, -21883, -24563, 
    -26373, -28316, -31159, -30107, -32007, -29151, -27446, -28031, -23363, 
    -22666, -17607, -16288, -12299, -7045, -2471, 2104, 5357, 9924, 13611, 
    18329, 21927, 24765, 26955, 28665, 30627, 30531, 30482, 31252, 27946, 
    27670, 24287, 21763, 18694, 14158, 9333, 7131, 2155, -2472, -6736, 
    -11334, -14011, -17805, -22540, -24898, -26235, -30523, -29499, -30304, 
    -30530, -31182, -29785, -25373, -23879, -21988, -19082, -14000, -13005, 
    -6984, -1928, 977, 6473, 10432, 14769, 17515, 20679, 24414, 26358, 28259, 
    30153, 31012, 30797, 31398, 29391, 27896, 24158, 21014, 20190, 16655, 
    10380, 7144, 2190, -2169, -6008, -10298, -14663, -17905, -22608, -24101, 
    -25972, -28693, -31053, -30238, -31787, -29790, -28631, -28795, -25860, 
    -21196, -20026, -14939, -11740, -7120, -4992, 1492, 4942, 10868, 14998, 
    17571, 22569, 23437, 26307, 29699, 30035, 29994, 31178, 31360, 29550, 
    29178, 24319, 23415, 17452, 15842, 12877, 7452, 2465, -63, -5879, -10621, 
    -14367, -16821, -21516, -24046, -25895, -28284, -29042, -31301, -30875, 
    -31138, -28410, -28827, -24706, -22347, -18023, -15086, -13119, -7878, 
    -3299, 1933, 5726, 10449, 12653, 17066, 20580, 25026, 26882, 26693, 
    29092, 31677, 30107, 30880, 29993, 26473, 26595, 22786, 19978, 16836, 
    11856, 7807, 4696, 114, -6375, -7878, -13048, -16488, -19608, -24170, 
    -24813, -28016, -28917, -29330, -31975, -30780, -28432, -27201, -26248, 
    -23218, -19759, -17511, -12641, -8331, -4533, 1010, 5018, 10216, 13721, 
    18143, 21390, 22516, 25941, 26959, 30711, 29906, 30997, 30319, 31138, 
    28665, 26902, 23029, 20188, 17763, 12348, 7593, 4309, -707, -5433, -8952, 
    -12429, -16622, -19651, -23344, -25181, -27323, -29938, -31493, -31626, 
    -30343, -29238, -28030, -25653, -23790, -19691, -17222, -12042, -8317, 
    -4755, -117, 4549, 7515, 11359, 15417, 19336, 21567, 26358, 27998, 28960, 
    30834, 30484, 30266, 28554, 29242, 25431, 24611, 21313, 15909, 12813, 
    8320, 3278, -31, -5259, -9632, -12448, -15376, -19106, -24172, -25115, 
    -26524, -30574, -30982, -31654, -29441, -29733, -27518, -25697, -23499, 
    -20011, -17631, -11822, -9085, -5969, -193, 3995, 7496, 11620, 15494, 
    18475, 22993, 25301, 29319, 29186, 30409, 31492, 30628, 30184, 28958, 
    26576, 24142, 20103, 17279, 13365, 7877, 4983, 723, -3633, -7640, -12013, 
    -16316, -20369, -22220, -26479, -27475, -30475, -30728, -31192, -29724, 
    -28692, -29445, -26358, -24807, -19998, -16366, -13940, -8610, -4965, 
    -704, 2641, 8852, 12011, 15168, 21114, 22599, 24373, 28636, 29276, 30244, 
    30567, 31192, 28334, 28868, 26757, 25148, 22083, 16497, 13778, 9834, 
    6616, 1848, -3181, -8393, -12229, -14489, -20139, -22949, -25910, -26929, 
    -29075, -30691, -30859, -31642, -28700, -28084, -26570, -23648, -21413, 
    -18806, -13376, -9042, -6011, -1431, 2493, 6571, 12629, 16088, 19755, 
    22178, 25683, 29220, 29554, 31613, 31916, 31711, 29537, 28707, 27003, 
    23083, 21351, 17054, 14897, 8949, 6679, 834, -1716, -7919, -10351, 
    -16030, -18681, -22206, -23888, -27886, -28547, -31197, -29651, -31701, 
    -30832, -30468, -26446, -23687, -22719, -17127, -13478, -9104, -6815, 
    -2314, 1179, 7803, 11260, 15593, 19649, 22558, 23558, 27346, 28615, 
    28966, 29870, 31481, 31403, 28659, 25625, 24839, 20685, 18024, 13733, 
    11155, 6153, 933, -2470, -7355, -11741, -15488, -17949, -22176, -26451, 
    -28091, -29473, -28968, -30082, -29920, -29864, -28624, -26113, -25795, 
    -21541, -18383, -14574, -12517, -6327, -3870, 1877, 6417, 11588, 14566, 
    18078, 20015, 24879, 26465, 28386, 30182, 31678, 30405, 30121, 28714, 
    27870, 25017, 22037, 19719, 13620, 12268, 5288, 1765, -1518, -6561, 
    -9269, -16408, -18205, -22564, -26066, -26524, -28950, -29190, -30216, 
    -29990, -29364, -28650, -26973, -23853, -21529, -18699, -14772, -11645, 
    -7230, -4194, 1361, 5685, 9551, 13139, 18183, 21672, 24275, 27558, 28971, 
    29664, 31218, 29533, 29400, 29458, 25978, 24457, 22342, 19155, 16408, 
    11172, 7695, 3047, -2879, -5985, -9827, -15454, -17116, -20038, -23778, 
    -26480, -28898, -30861, -31736, -32161, -30084, -29745, -27615, -24338, 
    -22190, -18728, -15085, -12444, -7226, -4225, 877, 5472, 10292, 13677, 
    18938, 21509, 23499, 26783, 28851, 29553, 30817, 29217, 29484, 28526, 
    29245, 24981, 24420, 18628, 16079, 10875, 8385, 3923, -1074, -7067, 
    -10817, -14245, -17069, -21745, -22696, -25529, -29292, -30129, -30982, 
    -30487, -30486, -28991, -27995, -25615, -22831, -20185, -15360, -11311, 
    -6383, -1854, 1008, 6450, 9658, 13568, 16332, 20618, 25077, 26234, 28480, 
    29369, 29550, 30628, 31246, 30129, 27538, 25579, 22097, 20209, 17185, 
    11288, 8558, 3784, -1096, -5365, -10159, -12232, -17455, -20469, -23907, 
    -25404, -29683, -29915, -29953, -30007, -31654, -30511, -28267, -24888, 
    -23077, -18961, -16505, -11272, -9116, -3984, -71, 4091, 10186, 13083, 
    17650, 21674, 23508, 24804, 27574, 30690, 32425, 30983, 30058, 30815, 
    28181, 25876, 23734, 19734, 15841, 11255, 6560, 2575, 15, -5551, -9002, 
    -11722, -17142, -20784, -24819, -24886, -27280, -30616, -30258, -31356, 
    -31020, -29850, -28097, -25670, -23901, -20118, -17372, -13420, -7224, 
    -6041, -1058, 3567, 9397, 13007, 16407, 21008, 23206, 26006, 27727, 
    29701, 29921, 31875, 30573, 29978, 28216, 25252, 22786, 19769, 17172, 
    13962, 9738, 4523, 1947, -3827, -7160, -13671, -15485, -19060, -23829, 
    -26756, -29158, -29063, -31476, -29474, -30173, -29912, -26462, -26286, 
    -23286, -20312, -16033, -14643, -10072, -5036, -247, 3071, 7035, 13758, 
    15382, 19608, 22893, 25930, 28728, 30629, 31480, 29634, 29918, 30193, 
    26983, 27281, 24226, 20689, 17299, 14388, 8894, 3878, 1080, -3891, -8739, 
    -12023, -15779, -18937, -21582, -23894, -28005, -27659, -29979, -30308, 
    -29582, -28281, -27777, -26347, -24054, -21814, -17328, -13616, -9153, 
    -5302, -660, 3829, 7941, 12043, 16128, 20042, 22853, 25938, 26341, 29555, 
    30474, 30462, 29542, 29252, 28507, 28146, 23866, 19057, 17863, 13472, 
    8601, 7096, 1597, -2284, -6886, -11860, -15587, -20066, -20768, -26633, 
    -28885, -30431, -29908, -31033, -29593, -28302, -29061, -25959, -24670, 
    -21737, -17642, -13418, -9242, -7247, -2086, 4142, 6944, 12616, 15761, 
    18992, 21964, 25449, 27048, 28808, 28938, 32054, 29110, 31195, 27852, 
    27889, 24091, 21056, 18690, 14298, 10400, 5943, 2820, -3381, -7878, 
    -11092, -15046, -19017, -22527, -24560, -27912, -29833, -29377, -29958, 
    -29997, -29286, -28973, -27337, -24158, -21210, -19253, -14869, -11429, 
    -6318, -1366, 2575, 6310, 12310, 14937, 18767, 22034, 23967, 27386, 
    29509, 30722, 29978, 29605, 29612, 28073, 27584, 25798, 20467, 17745, 
    13905, 11042, 6490, 3535, -1812, -7117, -11811, -15934, -18423, -23336, 
    -24571, -26387, -29014, -28538, -31053, -30078, -28871, -29551, -27203, 
    -25538, -21384, -18005, -14288, -12193, -6026, -2885, 2682, 7428, 10799, 
    15623, 18853, 21913, 26501, 25783, 29472, 30270, 29425, 30131, 31278, 
    29494, 27933, 25681, 22786, 18382, 14069, 9997, 7077, 1936, -2324, -6430, 
    -10733, -15411, -19140, -22102, -25287, -25979, -27658, -30345, -31492, 
    -29139, -29749, -28738, -27156, -26158, -23876, -18650, -15320, -10735, 
    -6220, -2346, 1655, 5912, 11161, 14486, 18681, 20854, 25164, 28114, 
    28380, 30073, 31182, 31995, 28792, 30124, 27427, 26630, 22224, 18600, 
    14079, 12533, 6889, 2894, -1221, -4633, -11520, -13824, -18707, -21904, 
    -25003, -26341, -27739, -30158, -31049, -29467, -31326, -28921, -27032, 
    -24054, -21925, -19593, -14025, -10976, -7380, -4054, 1810, 7591, 8304, 
    15237, 17933, 21388, 25022, 25538, 28580, 30408, 30747, 30644, 31011, 
    29535, 27734, 26264, 22927, 19267, 14698, 12943, 8226, 3299, -1368, 
    -6086, -8419, -13306, -18067, -20568, -24272, -25162, -28092, -29156, 
    -32259, -30055, -31587, -30419, -26539, -26747, -23158, -19499, -15583, 
    -12359, -7637, -3720, 2165, 5137, 9918, 13289, 16383, 21989, 24717, 
    26284, 29580, 28324, 30542, 30438, 30817, 28296, 27000, 24428, 22766, 
    20174, 15816, 12207, 6607, 4193, -446, -4454, -9269, -14908, -17140, 
    -21152, -23169, -26466, -27264, -28785, -31360, -30547, -29456, -29351, 
    -27357, -25527, -22311, -20488, -16476, -12813, -8017, -2845, -746, 4745, 
    8380, 12949, 17127, 20901, 21895, 26696, 27879, 29760, 30282, 31731, 
    30692, 30861, 28172, 26291, 23852, 19515, 17495, 13835, 7625, 4873, 
    -1079, -3898, -8461, -12315, -16663, -19616, -24851, -26088, -28773, 
    -29595, -29147, -31759, -31520, -29573, -27968, -24661, -23005, -20171, 
    -18255, -14149, -8502, -4130, -913, 3738, 8523, 13043, 17667, 19516, 
    22029, 26483, 27974, 30034, 30442, 29127, 30912, 30456, 27416, 25547, 
    25099, 20648, 16645, 13359, 10239, 4312, -73, -3806, -8965, -11338, 
    -16675, -20154, -22121, -24833, -29377, -30561, -30658, -30868, -32029, 
    -29850, -28673, -26375, -23108, -19715, -16545, -14328, -10374, -5478, 
    -489, 2667, 8280, 11499, 16074, 19396, 21484, 26020, 27618, 28887, 31366, 
    30618, 30816, 28474, 27309, 25991, 23987, 20854, 16815, 12631, 9057, 
    5979, 2436, -3456, -7923, -12948, -15463, -18005, -23352, -26576, -27259, 
    -28868, -29784, -30692, -30321, -29009, -29339, -26030, -23881, -20718, 
    -17711, -13817, -9336, -6084, -739, 5256, 6037, 11343, 16629, 18835, 
    23148, 25061, 27860, 29454, 29944, 31553, 31564, 30046, 28168, 27622, 
    23692, 21030, 18068, 14194, 9704, 6602, 1105, -3283, -7990, -12365, 
    -14828, -19656, -22519, -25194, -26800, -29942, -31302, -31960, -31218, 
    -29631, -27620, -25302, -24071, -20654, -17185, -14676, -10499, -5280, 
    -1226, 4293, 7527, 12675, 15592, 18634, 22406, 24907, 27041, 28985, 
    29403, 30861, 30629, 29429, 28623, 25866, 24163, 21257, 18028, 13205, 
    10685, 5851, 2468, -2733, -7789, -10246, -14191, -18837, -22215, -25018, 
    -26368, -28769, -30648, -29955, -32323, -30554, -29323, -28327, -24219, 
    -22381, -19049, -14274, -10818, -7686, -1439, 1959, 6945, 11869, 15586, 
    19648, 21810, 26158, 25975, 28516, 29172, 31260, 31331, 29877, 29561, 
    27816, 24395, 21736, 18270, 14165, 10008, 7744, 2670, -2495, -6442, 
    -10822, -14870, -17710, -22148, -24840, -27952, -28657, -31073, -31081, 
    -29300, -31544, -28171, -26696, -25600, -22774, -17263, -15056, -11156, 
    -7453, -2905, 2513, 6463, 10040, 14273, 17856, 21905, 24055, 26807, 
    30408, 29833, 31185, 30550, 29992, 27909, 27158, 24199, 23220, 18569, 
    14104, 11354, 7984, 1617, -1388, -6657, -10748, -15162, -19368, -21736, 
    -23797, -27864, -29372, -30212, -31045, -29386, -30663, -28809, -27674, 
    -25778, -21272, -18177, -15365, -11360, -7996, -2070, 586, 6101, 9345, 
    13899, 18416, 21316, 24711, 27512, 29537, 29784, 29845, 31162, 30965, 
    29315, 27207, 25492, 21144, 18432, 16386, 10283, 7977, 3073, -1512, 
    -6638, -9846, -15608, -16966, -21255, -25781, -25388, -29376, -28512, 
    -30448, -30430, -29905, -29475, -28492, -24368, -23089, -18836, -16278, 
    -11625, -7215, -3092, 2015, 6719, 10768, 14807, 18135, 20221, 23936, 
    25598, 29295, 29204, 31795, 30723, 29731, 29300, 28469, 25331, 22580, 
    20088, 16816, 11091, 7036, 4513, -270, -4132, -10656, -15020, -18284, 
    -21514, -22966, -26136, -28537, -30374, -31430, -31507, -29654, -28483, 
    -28061, -25371, -23452, -20757, -15339, -12445, -8478, -3919, -475, 4752, 
    9445, 14295, 16591, 19458, 24431, 27187, 29878, 29639, 29646, 29054, 
    31070, 28870, 27383, 24007, 21904, 19333, 16467, 12056, 7669, 4011, -379, 
    -4863, -8781, -12852, -18346, -20130, -24531, -26392, -29404, -30223, 
    -30916, -30407, -29454, -31201, -29441, -26433, -23451, -18905, -16334, 
    -13048, -6814, -4240, 349, 3943, 8953, 12788, 17058, 21081, 23351, 26429, 
    27754, 29237, 30976, 31493, 32006, 30217, 26232, 26815, 24551, 19213, 
    16536, 13533, 8740, 4693, -927, -4230, -8942, -12023, -17170, -19972, 
    -23650, -27152, -27270, -30167, -31832, -31344, -29279, -28342, -27260, 
    -26039, -23043, -20342, -18136, -12314, -8635, -4178, -993, 3266, 7908, 
    11693, 15287, 18728, 24667, 25262, 28255, 31055, 30357, 30252, 31007, 
    29998, 27034, 25920, 23654, 19895, 18538, 13900, 7835, 5077, -583, -4485, 
    -8530, -12534, -16677, -20559, -23298, -25290, -27967, -30939, -29552, 
    -29808, -31266, -29177, -26701, -25388, -24236, -20573, -15748, -12101, 
    -9196, -3505, -1878, 3823, 7445, 12774, 16961, 18581, 23791, 25474, 
    28520, 29556, 29464, 30011, 30840, 29616, 28812, 26415, 24771, 21653, 
    18193, 12796, 10956, 6462, 686, -3232, -8803, -11391, -16116, -19704, 
    -21720, -24659, -29211, -29140, -31860, -30957, -32243, -29146, -28003, 
    -26856, -23141, -21212, -17337, -13263, -9396, -5185, -2296, 3549, 8506, 
    11167, 15766, 19035, 22855, 26096, 27177, 29622, 31448, 32192, 29307, 
    29456, 28281, 27212, 23498, 21552, 16306, 13863, 10592, 6184, 1287, 
    -3806, -9123, -10786, -15751, -17560, -23652, -26289, -25730, -28591, 
    -30811, -31561, -30321, -30436, -26999, -27127, -23846, -20912, -17081, 
    -14135, -9755, -3903, -524, 3144, 6691, 11257, 15715, 19039, 22150, 
    26157, 27681, 28170, 30932, 30430, 30854, 30427, 27826, 26708, 25338, 
    21288, 17515, 13410, 9986, 5960, 3076, -2798, -7466, -11219, -15204, 
    -19212, -22872, -24933, -28516, -28828, -29518, -31589, -30051, -29996, 
    -27778, -26333, -23658, -20400, -19018, -13363, -8758, -6147, -952, 1756, 
    8000, 10961, 14083, 18176, 22767, 25009, 25651, 28310, 30716, 30811, 
    30481, 31122, 29375, 26014, 24280, 20958, 18812, 15787, 9951, 6124, 2330, 
    -1409, -7288, -10941, -16182, -18336, -20226, -23545, -28184, -29651, 
    -30506, -30731, -30561, -29422, -28659, -26049, -26011, -22139, -18625, 
    -13234, -11398, -6069, -1003, 1931, 7166, 10779, 14974, 18178, 20944, 
    24091, 26797, 27779, 30814, 30801, 30245, 30318, 27799, 25867, 23644, 
    22045, 17050, 15248, 10783, 7176, 1591, -3661, -5408, -11701, -14006, 
    -18247, -20752, -23008, -26846, -28369, -30442, -31237, -29732, -31729, 
    -28054, -27748, -24727, -22744, -17935, -15708, -11010, -8505, -3826, 
    447, 6323, 10733, 15186, 18166, 21398, 24343, 27443, 28227, 30592, 30757, 
    29949, 30944, 29080, 28914, 25341, 22146, 19810, 14243, 11723, 8868, 
    3562, -1506, -5678, -9448, -14915, -18471, -19646, -24011, -25747, 
    -27267, -28912, -31531, -30807, -30820, -28891, -27878, -25688, -21396, 
    -19740, -15064, -10445, -5806, -4227, 1996, 5962, 8727, 12901, 17140, 
    20999, 25056, 25647, 28505, 30410, 31317, 31008, 31897, 29140, 27856, 
    26444, 22831, 18888, 15962, 11882, 8839, 2545, -1238, -5885, -10763, 
    -13034, -17331, -19791, -23550, -27046, -29864, -29922, -30007, -30036, 
    -30608, -27970, -27009, -26216, -22925, -18419, -16267, -10701, -7657, 
    -2338, 1289, 5134, 10106, 13964, 17949, 21111, 24205, 26021, 29106, 
    28917, 30324, 30073, 31030, 29093, 28139, 26896, 23399, 19637, 16399, 
    10687, 8508, 2625, 157, -4620, -8989, -12517, -16985, -20626, -23624, 
    -26296, -27987, -28349, -29348, -32042, -31575, -29129, -27816, -26071, 
    -23889, -18428, -16942, -11697, -9165, -4146, 1586, 3106, 9503, 12409, 
    17156, 21957, 24102, 26570, 28358, 29566, 30918, 29686, 31544, 30587, 
    27365, 27044, 23856, 19305, 17296, 13665, 6849, 4254, 1232, -4714, -9407, 
    -13271, -17265, -21117, -22877, -24905, -28154, -27956, -31565, -30658, 
    -29487, -29683, -27717, -25295, -24403, -20276, -16993, -11587, -8037, 
    -3068, 1666, 4413, 7204, 13227, 15815, 20397, 22971, 24469, 27847, 29140, 
    31651, 30937, 30408, 28710, 29232, 26626, 23564, 19865, 17236, 12464, 
    9191, 3977, -705, -3570, -8278, -12688, -17795, -19307, -24310, -25545, 
    -27948, -30756, -31630, -31096, -30130, -28727, -29481, -24508, -22955, 
    -18616, -17084, -12402, -8631, -4784, -229, 4001, 9454, 13888, 16137, 
    18864, 21588, 25255, 27623, 29134, 29722, 31481, 31549, 29684, 29744, 
    27147, 23225, 20922, 17792, 13006, 10307, 5302, 961, -3406, -9276, 
    -11783, -16698, -20133, -22081, -26144, -27840, -28782, -30988, -31757, 
    -29562, -28156, -29012, -25674, -23388, -22211, -17575, -14489, -9006, 
    -3951, -960, 4897, 8862, 12525, 15734, 20212, 23592, 26258, 28723, 29149, 
    29555, 30824, 31351, 29192, 28228, 26009, 24494, 19909, 17527, 12602, 
    10032, 3848, 1061, -2559, -7395, -12064, -15623, -18482, -23781, -25983, 
    -27948, -29416, -30196, -31824, -29826, -30285, -28875, -25603, -22904, 
    -19964, -17981, -15371, -9839, -6124, -1158, 4346, 7072, 11797, 14993, 
    20150, 21720, 26761, 27398, 29507, 31455, 31276, 30888, 29098, 28147, 
    25689, 25195, 21520, 17176, 15443, 8963, 6968, -8, -2830, -8291, -10967, 
    -15539, -19621, -20718, -24553, -27244, -28707, -29826, -31529, -31824, 
    -30114, -28985, -27394, -23904, -21311, -18826, -14862, -10211, -5445, 
    -784, 2725, 7788, 12521, 16167, 20554, 22416, 24067, 26376, 29521, 29500, 
    32531, 30144, 30359, 29627, 26904, 23752, 23329, 18497, 14582, 11450, 
    6258, 3039, -3673, -5376, -9441, -14951, -19345, -20884, -24735, -27112, 
    -27924, -29898, -31009, -30637, -29466, -27508, -27140, -24920, -21255, 
    -20109, -14893, -9724, -5582, -2937, 2299, 7376, 10705, 14231, 18966, 
    21379, 24633, 26186, 29144, 30327, 29700, 31529, 29332, 29306, 27091, 
    23180, 22305, 18775, 14249, 10624, 7878, 1771, -2751, -5983, -10278, 
    -16401, -17605, -22148, -24841, -27640, -29244, -29800, -31543, -30743, 
    -30233, -28069, -26348, -23693, -22300, -20266, -15905, -11093, -8110, 
    -2604, 1587, 6363, 9657, 12498, 17070, 21353, 23607, 25729, 28190, 28661, 
    30257, 31169, 29147, 29386, 28157, 24815, 22778, 20357, 16674, 11767, 
    7965, 3497, -825, -5536, -11126, -13981, -17119, -20936, -24730, -26311, 
    -29963, -30647, -29546, -30640, -30046, -29964, -27368, -24640, -21855, 
    -19482, -15679, -11570, -7222, -3098, 897, 6838, 10217, 12500, 16984, 
    20320, 22767, 26226, 27024, 29019, 31652, 31158, 29214, 28732, 26207, 
    23551, 22560, 18351, 16217, 12494, 8386, 3889, 618, -4966, -9630, -14407, 
    -16587, -21381, -22698, -26941, -28850, -30346, -30436, -29327, -32036, 
    -28558, -27382, -25399, -23445, -19630, -14483, -12345, -8231, -3845, 
    -384, 5479, 8286, 15021, 17097, 20560, 22703, 26934, 26753, 29994, 29519, 
    29900, 31740, 29012, 28035, 23947, 21871, 20852, 16327, 11562, 6720, 
    3830, -667, -5284, -11013, -13862, -16109, -21643, -22563, -25726, 
    -27177, -28866, -31946, -31337, -29823, -29803, -28393, -25271, -23173, 
    -18833, -16824, -12874, -7690, -2243, 770, 5539, 9356, 12904, 17118, 
    19728, 24225, 26191, 28946, 31381, 29297, 29482, 32209, 28705, 28231, 
    24748, 24029, 20126, 14917, 13322, 9107, 4378, -454, -4605, -8921, 
    -14194, -17215, -22094, -23757, -25040, -28264, -30098, -29246, -30864, 
    -31852, -30233, -28292, -26353, -23836, -20154, -16182, -11539, -7051, 
    -3795, 1520, 5015, 7566, 12488, 16815, 18955, 23463, 25855, 29018, 29138, 
    30148, 30890, 30746, 28272, 28585, 26253, 23992, 19633, 16474, 14185, 
    9531, 5149, 1224, -5343, -7587, -12391, -17565, -20384, -23548, -26297, 
    -29765, -28675, -30311, -29422, -29856, -30479, -27937, -25443, -22346, 
    -19355, -15226, -14565, -9306, -3566, 632, 3767, 8989, 11830, 16226, 
    20737, 22016, 25565, 28586, 29323, 29768, 30675, 31360, 30976, 29763, 
    25533, 23609, 19785, 16453, 13877, 9470, 6090, 531, -4429, -9479, -11927, 
    -17808, -18650, -21715, -25271, -28079, -28337, -30935, -30669, -31942, 
    -29873, -29023, -25870, -24846, -20381, -17341, -14304, -10286, -7003, 
    -352, 4325, 7768, 11468, 15346, 20509, 23031, 26208, 27882, 28490, 30659, 
    30755, 30938, 29572, 28359, 26713, 23078, 20688, 16305, 12607, 9821, 
    4886, -531, -3434, -7332, -13220, -15299, -19556, -23742, -25367, -27137, 
    -29730, -31055, -29884, -30086, -29272, -28542, -26492, -23414, -20214, 
    -18680, -12753, -9880, -6532, -2248, 4441, 8427, 11090, 15324, 19106, 
    22892, 25136, 27416, 28572, 30374, 32178, 29203, 29487, 27054, 27432, 
    25513, 22453, 18571, 13560, 10137, 5529, 1484, -1694, -7752, -12322, 
    -15817, -18928, -21190, -26145, -28259, -30322, -30183, -31136, -30294, 
    -30498, -27319, -26708, -23821, -21439, -18153, -14403, -12088, -7242, 
    -2221, 2733, 6878, 11567, 15233, 19200, 21862, 24507, 27198, 29927, 
    28744, 30325, 30314, 28716, 28727, 26220, 23536, 23103, 17593, 15202, 
    11241, 6988, 2664, -1574, -6739, -9848, -14648, -20259, -21132, -25898, 
    -28234, -28695, -31091, -29969, -30794, -30433, -29340, -26154, -25166, 
    -21952, -18204, -15739, -9991, -8338, -1827, 1939, 5916, 10639, 14233, 
    17356, 22580, 25527, 27418, 27762, 28819, 31038, 30486, 30292, 28167, 
    27427, 26204, 21791, 16975, 14763, 11553, 4984, 1901, -622, -6481, 
    -10649, -13165, -18583, -21670, -24752, -25711, -27392, -30390, -31538, 
    -31795, -29207, -27945, -26802, -25253, -22670, -20250, -16569, -10106, 
    -6466, -3921, 1943, 6915, 11750, 13210, 18930, 22249, 24154, 26709, 
    29456, 31469, 29300, 30292, 30947, 30471, 26235, 25181, 23500, 19327, 
    15114, 12609, 6872, 2791, -1692, -5447, -10382, -14484, -17918, -20962, 
    -24334, -26065, -28464, -30953, -30372, -30182, -31084, -29438, -25844, 
    -24545, -22104, -18636, -16308, -10557, -7305, -4184, 2024, 4934, 10999, 
    14012, 17488, 19860, 23805, 25738, 28651, 29512, 32161, 30995, 30659, 
    28185, 28179, 24593, 23814, 19419, 15601, 12478, 9141, 3379, -245, -4501, 
    -9755, -13807, -18040, -20919, -24056, -27396, -29505, -29588, -29488, 
    -32200, -30305, -30537, -28493, -24735, -21148, -20381, -16580, -12783, 
    -6540, -2593, 710, 6639, 8878, 12351, 18456, 21038, 24259, 26432, 29364, 
    30496, 30620, 32311, 30052, 28445, 29284, 25662, 24295, 18220, 16022, 
    12268, 7438, 2916, 679, -5734, -9848, -12556, -17354, -19711, -23716, 
    -26367, -27959, -28484, -30847, -31637, -30444, -29367, -28227, -25887, 
    -22507, -20665, -16517, -12355, -8243, -3715, 941, 4990, 7920, 11613, 
    17571, 20953, 21733, 26833, 28832, 30437, 31297, 29691, 29270, 29141, 
    28786, 26420, 22115, 18976, 16206, 12435, 10014, 4249, 243, -4018, -9846, 
    -13550, -16189, -20323, -24626, -24589, -27832, -29679, -32109, -31247, 
    -29271, -29129, -28336, -25985, -24798, -19648, -16330, -13593, -8767, 
    -3859, 1162, 3981, 7914, 12840, 15770, 19848, 24019, 27125, 27043, 29778, 
    31235, 30552, 30227, 29550, 27758, 26776, 24464, 20841, 15124, 12488, 
    9851, 4052, -596, -4278, -9146, -12798, -16743, -20150, -23475, -25744, 
    -29421, -30004, -31674, -31613, -29355, -30624, -27023, -26821, -22958, 
    -20335, -17486, -13588, -8335, -5968, -477, 2080, 6464, 12028, 16127, 
    20553, 22375, 25463, 28041, 29485, 29147, 31149, 30610, 28840, 29163, 
    25301, 23605, 19804, 17279, 12173, 8807, 3959, 1970, -2364, -8012, 
    -13147, -17656, -20519, -22207, -25426, -27302, -28166, -30290, -32178, 
    -29753, -31083, -28265, -26741, -24695, -21077, -17510, -13888, -9502, 
    -3845, -456, 4312, 6851, 10511, 16366, 19703, 23195, 24962, 27126, 30497, 
    30364, 29900, 31010, 29902, 29690, 27199, 23911, 20792, 17235, 14091, 
    10137, 5663, 1551, -3309, -8720, -11218, -14904, -19200, -22844, -24788, 
    -26265, -30391, -29285, -30790, -31733, -29322, -27886, -25560, -24642, 
    -22179, -18918, -13282, -10275, -5782, -2186, 2800, 7889, 11283, 16499, 
    19822, 22801, 24672, 26710, 28829, 29893, 30488, 29887, 31058, 28571, 
    26533, 25680, 22072, 16697, 14175, 8633, 5513, 1061, -3158, -7454, 
    -12005, -14846, -18958, -22792, -25258, -26689, -29329, -31226, -31529, 
    -31437, -29416, -27337, -28000, -23736, -21342, -19171, -14629, -9390, 
    -6179, -1617, 3425, 6933, 10935, 14267, 17643, 22604, 25606, 28390, 
    29606, 29985, 30895, 29719, 28918, 28136, 26830, 23970, 20554, 17781, 
    13068, 11330, 6140, 2608, -2373, -8085, -10968, -14709, -17155, -22305, 
    -23704, -25906, -28150, -29384, -29698, -30474, -31281, -28503, -26247, 
    -23790, -21227, -18613, -14701, -12055, -6232, -2457, 1493, 6254, 10532, 
    15671, 19093, 22357, 24613, 26445, 29552, 30021, 31360, 31018, 30487, 
    28064, 26205, 24491, 22442, 19700, 13407, 11115, 6211, 2697, -287, -7275, 
    -9614, -14658, -19146, -22692, -23671, -27849, -28198, -30743, -30309, 
    -31491, -29505, -29023, -27699, -24494, -21967, -19190, -13959, -12881, 
    -7913, -2743, 1622, 7299, 10475, 13912, 18871, 20726, 25276, 28105, 
    30036, 31431, 30213, 29710, 31744, 28860, 27295, 23987, 22278, 18827, 
    16609, 10351, 7178, 2518, -1717, -5337, -10199, -14810, -17204, -21161, 
    -25706, -25965, -28801, -30903, -32127, -30303, -30149, -27801, -28755, 
    -26757, -21956, -19750, -15125, -12312, -8424, -3255, 184, 4439, 10701, 
    12538, 16412, 21193, 23032, 26630, 28289, 30487, 30873, 31566, 30709, 
    29014, 27234, 25137, 22347, 19957, 15308, 11022, 7886, 4133, -725, -5900, 
    -10919, -12725, -18491, -21654, -23995, -25499, -27550, -30283, -31568, 
    -31860, -31120, -29054, -28003, -24839, -22985, -19614, -16441, -12195, 
    -8747, -2836, 336, 5467, 8435, 13142, 15859, 21941, 24823, 26428, 27568, 
    30041, 30867, 31134, 30315, 29455, 28550, 25699, 22422, 19852, 16377, 
    12100, 8424, 2286, -1806, -4436, -9350, -14993, -17172, -20941, -22940, 
    -27373, -28860, -29418, -31036, -31719, -32177, -29366, -28188, -26210, 
    -24218, -20685, -17042, -11791, -9074, -3902, 1279, 2985, 9099, 14216, 
    17747, 20766, 23526, 26850, 29333, 31345, 31748, 31002, 29131, 29728, 
    28181, 24658, 24574, 19476, 14894, 12327, 9590, 4891, -740, -4449, 
    -10271, -12376, -17539, -20437, -23099, -24237, -27716, -30599, -30196, 
    -31006, -29875, -30489, -28990, -27172, -22474, -20335, -17014, -12096, 
    -8602, -2883, -1293, 5599, 7541, 13409, 16041, 19549, 24399, 24931, 
    28824, 29258, 31033, 29496, 31037, 29539, 29345, 25948, 21961, 20174, 
    16204, 12453, 9923, 4445, -908, -5014, -8708, -11802, -16801, -21030, 
    -23190, -26127, -28940, -28314, -31384, -30533, -30479, -29295, -28018, 
    -25909, -22729, -20304, -17928, -12843, -9725, -4494, 290, 2513, 9620, 
    13203, 16086, 20426, 22432, 25439, 29596, 30309, 31143, 31189, 31082, 
    29802, 27635, 26135, 24037, 19380, 16676, 13133, 10040, 5306, -949, 
    -4338, -6492, -12479, -17535, -20326, -22561, -26395, -26081, -29333, 
    -29927, -31191, -32293, -31564, -28162, -28229, -23822, -20563, -16067, 
    -11928, -9074, -5368, -2039, 3444, 8596, 12475, 17038, 19561, 21986, 
    25148, 28416, 29448, 30371, 29735, 30018, 31246, 27738, 24942, 22989, 
    19439, 17029, 14286, 8696, 5796, 1537, -3820, -7937, -11656, -15323, 
    -18172, -22198, -26398, -27458, -30529, -30214, -30972, -29812, -29304, 
    -27920, -26613, -24091, -19470, -17552, -15074, -8506, -5406, -2033, 
    4214, 7671, 11193, 15253, 19847, 20958, 25795, 26866, 29068, 30854, 
    29084, 30856, 30619, 28580, 25564, 23811, 22332, 17660, 13935, 10037, 
    5072, 3, -2875, -6278, -12796, -14121, -18753, -22360, -25714, -26330, 
    -28280, -29244, -30223, -30061, -29101, -27744, -26358, -25545, -22213, 
    -16998, -14839, -9067, -6003, -1989, 4303, 7083, 10740, 14909, 19812, 
    21664, 25172, 26937, 28391, 30505, 29220, 31038, 29988, 29335, 26733, 
    23369, 21990, 19332, 14373, 10903, 5641, 1483, -2014, -7525, -10934, 
    -14867, -17655, -20663, -24493, -27900, -28351, -31712, -29645, -30531, 
    -30421, -29131, -27542, -24921, -22489, -17480, -14845, -9347, -6805, 
    -3091, 2560, 6223, 11788, 14847, 19518, 21806, 25210, 28056, 29869, 
    30022, 30850, 31641, 30006, 29160, 27889, 25902, 21362, 19486, 14212, 
    11011, 5662, 2027, -2524, -6216, -11542, -14334, -18535, -20392, -24355, 
    -26289, -29044, -30627, -30684, -30633, -29670, -30290, -26875, -26613, 
    -21647, -17957, -15620, -12078, -6859, -2053, 197, 5312, 9780, 14363, 
    18221, 20496, 24037, 27545, 27590, 29680, 31843, 30498, 30490, 30288, 
    26105, 24999, 21811, 19724, 15516, 10942, 6293, 2437, -2742, -6358, 
    -11029, -14137, -17274, -21807, -23932, -26686, -28189, -31171, -30613, 
    -30056, -30557, -28129, -27833, -24973, -21064, -18647, -16449, -11785, 
    -6228, -3787, 1342, 6556, 11263, 12663, 17341, 21857, 23111, 26386, 
    28251, 31467, 30946, 32393, 30485, 29005, 26116, 25900, 21728, 19206, 
    14871, 11625, 6931, 4092, -670, -5915, -8799, -14735, -17670, -21693, 
    -24638, -27171, -28640, -30328, -29727, -31475, -31626, -28503, -27956, 
    -25983, -22804, -19142, -15794, -12102, -8107, -3483, 1457, 5125, 8949, 
    13692, 17164, 20657, 24131, 26755, 28881, 29081, 31013, 31492, 29796, 
    29447, 28496, 24572, 22440, 19216, 15384, 13312, 7705, 4293, -924, -5122, 
    -8154, -13754, -16562, -21183, -25234, -26291, -28727, -30058, -31290, 
    -32099, -29839, -27800, -27992, -24706, -22981, -18929, -16078, -12423, 
    -7809, -4146, 540, 4884, 8766, 12961, 16890, 20458, 23517, 27118, 27122, 
    30487, 32048, 30269, 30044, 29709, 29001, 27072, 23913, 19479, 16778, 
    12140, 7610, 2759, -820, -5560, -7959, -14545, -16618, -20464, -22730, 
    -25297, -28743, -29560, -30256, -31244, -30443, -29997, -27947, -25983, 
    -23100, -20360, -17282, -12589, -9462, -5449, 276, 4507, 7806, 13041, 
    16184, 20228, 23923, 26554, 29076, 29430, 31515, 30704, 31337, 30784, 
    27156, 25725, 23858, 21753, 16705, 11734, 7981, 3796, -268, -3877, -8395, 
    -13834, -16303, -19783, -23486, -25032, -28194, -29701, -31683, -30629, 
    -30140, -29196, -27477, -24800, -24394, -20431, -16889, -14145, -8186, 
    -4779, -1230, 4481, 8754, 13336, 16227, 17937, 23845, 26667, 27522, 
    28970, 30001, 30837, 32349, 29484, 28504, 25294, 22172, 19344, 17356, 
    14909, 9664, 4323, 1492, -3499, -9421, -11249, -15880, -19023, -21754, 
    -25237, -27424, -28182, -28772, -29312, -29891, -29610, -26803, -27949, 
    -22654, -20547, -16096, -14297, -9706, -6488, -1598, 3889, 6593, 10989, 
    16369, 19494, 24274, 25200, 28231, 29526, 30566, 30553, 31837, 30283, 
    28901, 25935, 22967, 21104, 18037, 12936, 9675, 6717, 833, -3501, -7792, 
    -11552, -16109, -19673, -21469, -26307, -27776, -28845, -31958, -30779, 
    -30697, -29084, -28085, -25666, -24903, -21225, -16850, -13994, -9622, 
    -6402, -423, 2572, 7873, 11047, 16175, 18056, 21228, 26701, 27190, 28100, 
    29835, 31054, 29722, 29487, 27472, 27038, 24438, 22478, 16914, 13194, 
    11013, 5881, 1731, -3514, -6208, -11797, -13567, -19543, -23538, -25694, 
    -28370, -30030, -30439, -29148, -29894, -30303, -29508, -25909, -23819, 
    -21166, -19330, -14801, -10094, -5959, -2096, 2757, 6739, 10876, 14997, 
    17547, 23086, 25458, 26242, 28678, 29966, 29951, 29556, 30016, 29342, 
    26698, 23800, 20771, 18152, 13843, 10570, 6939, 1999, -1336, -7409, 
    -10380, -13925, -19611, -21395, -24504, -27233, -29012, -30007, -28897, 
    -29569, -31137, -29591, -26968, -25110, -22643, -17980, -16276, -11751, 
    -7394, -1659, 2478, 7109, 11273, 14972, 18762, 22724, 24897, 26843, 
    28830, 30719, 31426, 30853, 28464, 28479, 26525, 23677, 20192, 19112, 
    14977, 11853, 5515, 2346, -2697, -6812, -10717, -14630, -17742, -20354, 
    -24874, -26814, -28839, -31103, -32019, -31872, -30995, -28077, -27468, 
    -26792, -21835, -17480, -13834, -11914, -5514, -2210, 2074, 7445, 9635, 
    13807, 18604, 21633, 23441, 27220, 27190, 28798, 30633, 30608, 30866, 
    28897, 28202, 24405, 22829, 18445, 15645, 11933, 6385, 1351, -2349, 
    -7008, -9880, -15269, -18462, -22476, -23945, -26372, -28179, -30687, 
    -31526, -30928, -29899, -29257, -29077, -24207, -22954, -20024, -16523, 
    -13024, -7202, -3651, 2443, 6424, 10100, 14578, 16575, 20531, 25152, 
    26814, 28505, 28379, 30662, 30180, 31013, 30408, 27603, 25565, 23011, 
    17867, 16240, 11243, 6679, 3564, -651, -5546, -9077, -12880, -17930, 
    -21635, -25812, -26524, -27191, -30420, -30665, -30482, -29983, -28292, 
    -26118, -25255, -21784, -18939, -16701, -12121, -8604, -3583, 881, 4226, 
    9919, 13648, 16943, 21140, 24633, 26370, 28789, 29755, 31803, 31964, 
    31071, 29415, 27867, 27034, 22571, 19555, 16519, 13165, 7728, 3783, 
    -1162, -4566, -9101, -13299, -16637, -20439, -24804, -26488, -28064, 
    -27840, -31570, -30964, -29720, -29114, -26745, -25301, -22716, -18029, 
    -14624, -12177, -7812, -4536, 1949, 5273, 8621, 13392, 16775, 19690, 
    24462, 25567, 29103, 29191, 30042, 29755, 30585, 28956, 28664, 25656, 
    22291, 19195, 15055, 13427, 7018, 5830, -979, -3445, -10108, -13830, 
    -16994, -20454, -24237, -25716, -28250, -29412, -30188, -30616, -30275, 
    -29778, -27967, -25311, -23259, -20348, -16292, -12561, -8324, -4137, 
    680, 3010, 8949, 11080, 16830, 19402, 23008, 26025, 29453, 29906, 30624, 
    31649, 30584, 28815, 28590, 26982, 22597, 19888, 16006, 12303, 9055, 
    5879, 945, -3571, -8046, -11669, -17569, -18704, -24557, -26003, -27809, 
    -31013, -31152, -31008, -30687, -29662, -28075, -25225, -24281, -21292, 
    -18214, -11627, -9355, -5285, 259, 3061, 7586, 12574, 16412, 19129, 
    23125, 26024, 28003, 29291, 31964, 31957, 29394, 30707, 28988, 25425, 
    23742, 20335, 15948, 14718, 10519, 4432, 877, -3893, -9004, -10879, 
    -17499, -20249, -23624, -24357, -27505, -30000, -30088, -31380, -31330, 
    -29405, -27916, -27518, -23261, -21671, -17869, -13673, -8323, -5348, 
    -1870, 3129, 8702, 10523, 15506, 19033, 20939, 26417, 27607, 28946, 
    30474, 31176, 29634, 29353, 29538, 26679, 23588, 20006, 17431, 12319, 
    10167, 6144, 417, -2801, -7179, -10415, -15556, -18176, -23327, -25806, 
    -29335, -28050, -29453, -31221, -30062, -29365, -28746, -25712, -23548, 
    -21778, -16931, -15041, -9635, -5334, -1167, 3534, 7887, 12634, 14498, 
    19921, 21342, 24386, 28206, 28670, 30709, 30258, 31138, 30306, 29199, 
    26910, 24599, 21887, 18736, 13698, 8555, 5566, 2591, -2408, -7977, 
    -10106, -15553, -18787, -21115, -25591, -27833, -28664, -29592, -31430, 
    -30528, -30517, -28627, -26400, -24717, -21817, -19128, -13981, -10644, 
    -5932, -862, 1686, 6678, 11132, 15335, 18233, 21917, 24213, 26565, 29700, 
    29776, 32132, 31136, 30332, 28562, 26440, 24799, 21152, 18677, 13841, 
    11136, 7402, 1603, -1686, -6941, -11322, -14714, -18702, -23410, -24876, 
    -27119, -29304, -29999, -30090, -29583, -30007, -29038, -27070, -23070, 
    -22787, -18853, -15198, -9468, -5973, -2046, 1647, 5221, 10040, 16384, 
    18003, 21642, 26173, 27137, 29698, 30417, 31091, 29818, 30375, 29835, 
    25433, 23815, 20526, 19001, 15591, 11472, 7368, 3182, -1721, -6060, 
    -10330, -13926, -17395, -20626, -25569, -27346, -29585, -31066, -30427, 
    -30444, -28847, -28358, -27447, -26280, -23982, -19451, -15446, -11356, 
    -7205, -2014, 1818, 6116, 9232, 14573, 17109, 21317, 24672, 25282, 28880, 
    30257, 30851, 29531, 30527, 28512, 26913, 24522, 23812, 18499, 15636, 
    10843, 5649, 3657, -1759, -5322, -9646, -12935, -16650, -20993, -23694, 
    -27166, -30225, -30471, -29792, -31087, -30381, -29448, -27707, -25736, 
    -22916, -18915, -14869, -12204, -7919, -2808, 1562, 6111, 11300, 12871, 
    16317, 19650, 25324, 26869, 27917, 30033, 31015, 29663, 30343, 29869, 
    27578, 26442, 23092, 18309, 17207, 12149, 8178, 1568, -1558, -6394, 
    -8472, -13781, -18528, -20709, -24608, -26695, -28594, -29806, -30508, 
    -30595, -31460, -30208, -27198, -25734, -23505, -19415, -15217, -11730, 
    -6747, -2767, 1531, 6752, 10462, 13687, 18160, 20487, 24629, 26632, 
    29226, 29654, 30553, 32641, 30624, 28010, 27617, 26427, 22359, 18956, 
    17045, 13288, 8011, 2965, -337, -5145, -9189, -13075, -16074, -19296, 
    -23748, -25125, -28365, -29982, -31807, -30191, -29669, -30204, -29463, 
    -24582, -23358, -19805, -16622, -13512, -6958, -4102, 1560, 3144, 8187, 
    11787, 17527, 22078, 24126, 24877, 28055, 29618, 30795, 30062, 28870, 
    29153, 28342, 24681, 21810, 18848, 15190, 11745, 7027, 4836, -108, -4078, 
    -8774, -14194, -17519, -19890, -22817, -24672, -28248, -29105, -29959, 
    -30836, -31006, -29966, -28310, -27272, -22932, -20295, -16788, -11917, 
    -7644, -5399, 5, 3364, 8889, 11956, 17045, 21408, 24652, 26220, 28349, 
    29985, 30164, 31061, 31753, 29713, 27420, 26425, 23025, 20063, 16514, 
    12542, 7977, 5280, 237, -3871, -8200, -12743, -16576, -20297, -23160, 
    -25254, -26782, -28590, -30614, -31353, -30865, -28850, -27421, -25614, 
    -23516, -21756, -16507, -14503, -8986, -4364, -1564, 4590, 9321, 13205, 
    16724, 19981, 23975, 26188, 28975, 28882, 30073, 29952, 32110, 28896, 
    29134, 25568, 23932, 21985, 18171, 12416, 9956, 5394, 634, -3180, -8715, 
    -11667, -15682, -20080, -21555, -25525, -27609, -30047, -30498, -30884, 
    -30490, -29222, -29339, -27418, -23750, -21648, -17871, -14356, -10231, 
    -4879, 17, 3751, 6913, 11837, 16677, 19402, 23687, 26471, 28913, 28298, 
    30641, 29747, 30151, 31074, 26978, 26773, 23020, 20283, 17921, 14592, 
    11141, 4853, 877, -2819, -8611, -11585, -16697, -20364, -22038, -24372, 
    -27724, -28767, -28746, -29911, -30564, -29452, -26897, -27892, -24412, 
    -20126, -17163, -13475, -10102, -7115, -2320, 3805, 5670, 11881, 15522, 
    18411, 23920, 24436, 28044, 29638, 31727, 32165, 30873, 28260, 28520, 
    26211, 23064, 20964, 18108, 13913, 9118, 6729, 1197, -2642, -6301, 
    -11307, -15959, -20242, -22954, -24846, -27608, -29072, -29028, -31764, 
    -31143, -31007, -30100, -28136, -23965, -20824, -19605, -13569, -11592, 
    -5865, -3217, 2012, 6055, 11674, 14090, 19166, 21491, 25467, 27481, 
    28845, 29617, 31002, 31245, 28720, 29219, 26832, 24623, 22832, 19398, 
    14528, 10426, 6267, 2328, -2804, -7777, -10809, -15388, -19486, -21984, 
    -24986, -28245, -29066, -30472, -31005, -30129, -30477, -29368, -26932, 
    -24312, -20446, -19581, -13199, -9724, -6863, -3506, 3033, 6024, 11341, 
    14771, 17461, 23095, 25671, 25504, 30430, 28758, 30331, 30263, 30690, 
    28558, 25918, 24924, 22787, 17969, 14060, 10478, 6395, 1213, -1626, 
    -5402, -10783, -14640, -17865, -21654, -24649, -26660, -27220, -28807, 
    -31443, -29982, -29584, -29231, -26628, -25381, -22185, -18319, -15106, 
    -10923, -6677, -2129, 403, 7431, 10084, 14549, 19710, 23017, 23253, 
    26641, 29940, 29679, 29134, 30710, 30597, 28159, 27443, 23993, 22575, 
    19646, 16438, 11839, 7460, 1770, -1703, -7708, -8805, -15397, -18844, 
    -21723, -25090, -27513, -27540, -29651, -31621, -31337, -30123, -28084, 
    -27825, -26016, -22396, -18699, -16541, -12041, -8049, -4070, 2238, 4432, 
    10752, 15036, 18584, 21200, 23570, 26907, 28979, 30046, 30741, 30737, 
    30780, 27499, 28644, 26444, 21471, 20566, 15082, 12911, 8167, 3797, -971, 
    -5556, -9570, -14492, -16249, -21798, -23154, -26010, -29634, -29242, 
    -30176, -30981, -29391, -29532, -26515, -25355, -23037, -20576, -15627, 
    -10976, -6589, -3522, 107, 4465, 8378, 12588, 16792, 21381, 24271, 27739, 
    28345, 31056, 30383, 30495, 29248, 28837, 27528, 25272, 23992, 20360, 
    16427, 13571, 7960, 3036, -1738, -4857, -8435, -13073, -18382, -20504, 
    -23498, -26302, -29019, -30631, -29811, -30038, -29716, -28960, -27250, 
    -26649, -23208, -20439, -16264, -11930, -7084, -4461, 1522, 4016, 9317, 
    13203, 17304, 20943, 23258, 26107, 26548, 29734, 29496, 30518, 30315, 
    30000, 27914, 24035, 23819, 21261, 16310, 12592, 8919, 4380, -766, -5362, 
    -8451, -12620, -18177, -21015, -22086, -27309, -27590, -29289, -30016, 
    -30982, -30962, -29722, -27630, -24063, -22844, -19376, -16022, -13686, 
    -9222, -4769, 1731, 4752, 7158, 11938, 16994, 19757, 22295, 25517, 27523, 
    28240, 30074, 29602, 29505, 28351, 28459, 27461, 24172, 20896, 16690, 
    12323, 9393, 5418, 710, -3258, -8772, -11486, -16322, -19553, -23259, 
    -24586, -29072, -30265, -30050, -31239, -31302, -30674, -28552, -24956, 
    -23002, -19821, -17863, -11957, -9334, -4191, -316, 3858, 6733, 10733, 
    15355, 18789, 24286, 27116, 28439, 29088, 30499, 29986, 30983, 30102, 
    28694, 25728, 22685, 22063, 16610, 13182, 8824, 4787, 131, -3956, -7097, 
    -11617, -17669, -19644, -22291, -26293, -27155, -30867, -30440, -30884, 
    -30432, -29757, -27468, -25983, -22747, -20876, -17042, -13872, -8455, 
    -4974, -1998, 3347, 8753, 12402, 14911, 18238, 22299, 26100, 28408, 
    27943, 30600, 30390, 29545, 29964, 28721, 26855, 24972, 20688, 16288, 
    15438, 8177, 6113, 2019, -4298, -8499, -12165, -14505, -19657, -21448, 
    -24919, -27146, -29087, -31076, -31116, -31306, -29987, -29586, -26643, 
    -24304, -19923, -17697, -14120, -11158, -5240, -1437, 3354, 7589, 12210, 
    15359, 19064, 21134, 25169, 26971, 29225, 30387, 30207, 30973, 31168, 
    28448, 26400, 24668, 22388, 18764, 14662, 9906, 5958, 719, -2438, -7460, 
    -11338, -15035, -18303, -21316, -23954, -27331, -28634, -29808, -31253, 
    -30716, -30379, -28492, -25786, -23138, -22524, -18796, -14278, -11266, 
    -6437, -473, 2672, 6040, 10343, 14981, 18215, 21502, 26095, 27951, 30168, 
    30250, 31294, 31090, 29971, 30215, 27234, 23773, 21685, 19409, 14197, 
    9628, 4577, 1480, -2369, -5430, -10722, -15966, -18715, -22280, -24185, 
    -27996, -28887, -29291, -32075, -29778, -29046, -30002, -26402, -23793, 
    -21675, -20004, -15473, -9139, -7682, -2270, 2724, 8236, 10275, 15453, 
    18893, 23122, 24695, 27246, 29634, 30676, 29537, 31284, 28870, 29274, 
    25746, 25340, 21494, 18280, 15760, 10681, 6487, 2187, -1472, -5519, 
    -12269, -14457, -19350, -22638, -24121, -27344, -28953, -30716, -31841, 
    -29364, -30649, -27913, -27290, -25114, -22288, -18344, -15375, -11974, 
    -6401, -3593, 1338, 6245, 10835, 14513, 18980, 21525, 24752, 27376, 
    28678, 29523, 31204, 30174, 29856, 29040, 28702, 23690, 21063, 20301, 
    15387, 12883, 6923, 3761, -1851, -7683, -9976, -14727, -17102, -23021, 
    -24774, -27615, -28327, -29954, -30610, -29904, -31012, -28825, -26857, 
    -25405, -23367, -18911, -15418, -11250, -7256, -1162, 1541, 5040, 9436, 
    13682, 18394, 21854, 24250, 26247, 28679, 28537, 31884, 30393, 31109, 
    28673, 26827, 25276, 22851, 19442, 14439, 12492, 6994, 2592, -783, -4398, 
    -9232, -13767, -18620, -21575, -23256, -26148, -28019, -29775, -31106, 
    -31674, -31379, -28870, -27428, -26105, -22070, -20853, -16828, -13141, 
    -6271, -4342, 481, 6179, 8710, 13865, 16259, 21089, 24436, 24892, 28987, 
    29666, 29933, 31234, 30943, 29574, 28169, 24338, 23370, 19308, 16526, 
    11391, 6946, 3838, -1093, -5975, -9748, -12803, -17172, -21287, -24377, 
    -26345, -28305, -29181, -30419, -29743, -31788, -29788, -28360, -26258, 
    -22124, -21279, -17159, -11111, -8488, -3603, 1155, 6546, 9059, 14309, 
    17289, 20867, 22843, 24991, 27969, 30878, 29699, 30563, 29350, 29764, 
    26832, 26654, 22972, 20233, 16153, 12197, 8671, 5118, -627, -4160, -8384, 
    -13698, -18547, -20334, -23557, -25835, -28873, -30750, -29610, -30777, 
    -30741, -30233, -27427, -25219, -23316, -19693, -17003, -13411, -7251, 
    -5535, 345, 4374, 8480, 13060, 18257, 20401, 23341, 25902, 29400, 29279, 
    30667, 32053, 30993, 29420, 27601, 26197, 23512, 19467, 18006, 12846, 
    8004, 4962, 294, -4250, -8317, -11948, -16942, -20373, -23270, -24509, 
    -27559, -30964, -30260, -31463, -31209, -29204, -28511, -25870, -23111, 
    -20949, -17501, -12761, -8651, -4249, -632, 4797, 7746, 12747, 15375, 
    20558, 22356, 27065, 28942, 29565, 31668, 30563, 32150, 30101, 29234, 
    25961, 23549, 20610, 16844, 12397, 9874, 4955, 652, -3269, -9235, -11552, 
    -16014, -19782, -22771, -25320, -27296, -28510, -31468, -30465, -31563, 
    -29993, -28421, -26641, -24598, -19264, -18309, -14813, -9849, -3756, 
    766, 3514, 7325, 12266, 15039, 19689, 21819, 24045, 27332, 28683, 30716, 
    30069, 30524, 29601, 26744, 25292, 22803, 21172, 17755, 14384, 9894, 
    5559, 1956, -3625, -5818, -11213, -15440, -21005, -21893, -25803, -28031, 
    -29190, -29292, -31137, -30602, -29055, -29438, -25687, -23527, -19636, 
    -18022, -12693, -10886, -5873, -1338, 3035, 7699, 11605, 16913, 18678, 
    22206, 25513, 27545, 29127, 30171, 30024, 30655, 29925, 28718, 26150, 
    24175, 21034, 17033, 14136, 10502, 7278, 3222, -1982, -8057, -10447, 
    -15471, -18925, -21478, -25671, -26886, -29927, -30273, -29173, -31121, 
    -30617, -29042, -27492, -23070, -20900, -18946, -14493, -11458, -6384, 
    -2221, 3148, 7255, 12277, 15944, 17745, 22850, 25006, 27576, 28466, 
    29786, 30643, 29412, 31164, 27498, 27252, 23612, 20704, 19496, 14757, 
    9340, 7467, 1295, -1927, -5712, -10366, -14166, -18901, -22304, -25153, 
    -28538, -28534, -30474, -31858, -30362, -28763, -27605, -26640, -25706, 
    -22554, -18764, -14901, -10113, -7218, -2997, 2579, 7451, 11446, 13611, 
    18584, 21773, 24699, 26359, 29735, 28958, 29947, 30182, 28779, 29162, 
    27399, 24769, 21020, 20359, 13491, 10539, 8292, 2338, -1877, -5165, 
    -9098, -14855, -18334, -20659, -25762, -26910, -28126, -29978, -31134, 
    -30378, -30784, -28804, -27056, -25636, -22392, -20184, -15890, -11696, 
    -5828, -2290, 2116, 5863, 11116, 15092, 18245, 20871, 23688, 27229, 
    29971, 30457, 31983, 31258, 29832, 30500, 26436, 24014, 22385, 19621, 
    16734, 12134, 6725, 3694, -2900, -4567, -9383, -12706, -17901, -21856, 
    -23788, -26239, -28427, -30375, -31596, -29463, -30518, -28859, -28673, 
    -24970, -22378, -19680, -16800, -11977, -6393, -3920, 1379, 6209, 9335, 
    14269, 18072, 20879, 23301, 27321, 27700, 30048, 31225, 31280, 29868, 
    30521, 27605, 26061, 23502, 18519, 15684, 10536, 7382, 4402, -1468, 
    -4440, -11061, -12859, -17702, -21213, -23702, -27639, -27263, -30807, 
    -32302, -31544, -30728, -29567, -28230, -25155, -23336, -20054, -16582, 
    -11912, -8210, -1778, 986, 4592, 10355, 13244, 16624, 21704, 24125, 
    25903, 27997, 28960, 31479, 30270, 30105, 29795, 27798, 26060, 21575, 
    21287, 15950, 12251, 7651, 3573, -193, -5186, -9928, -14087, -15862, 
    -20495, -22905, -25859, -28397, -30325, -30482, -30805, -31015, -30462, 
    -26352, -24704, -22092, -20156, -16511, -12935, -8168, -4037, 310, 4372, 
    9039, 12219, 17634, 20291, 22568, 24444, 27617, 30319, 29316, 30200, 
    28893, 29313, 28688, 26192, 21728, 18966, 16115, 14046, 9552, 4113, 388, 
    -3113, -8692, -14296, -17312, -19579, -22201, -25983, -28435, -30716, 
    -29582, -29823, -29806, -31166, -29289, -25205, -22690, -18691, -15600, 
    -12769, -9540, -3430, -1351, 5332, 9764, 12466, 16119, 19712, 24418, 
    26209, 28794, 29259, 32007, 31186, 30177, 28866, 27930, 26531, 22640, 
    21298, 16928, 11766, 9729, 4296, -182, -4461, -9021, -12637, -17797, 
    -20268, -23194, -25603, -27581, -30124, -30330, -31005, -30701, -30331, 
    -27835, -26139, -24777, -20466, -16261, -13363, -7937, -6349, -205, 3992, 
    7911, 13026, 17050, 20240, 22927, 25655, 27295, 29763, 30263, 29120, 
    30079, 28818, 29322, 27035, 23048, 20125, 16399, 14498, 8401, 6339, 1089, 
    -2957, -7927, -12105, -17539, -20863, -22240, -26665, -27245, -28793, 
    -30055, -30421, -29906, -28976, -27253, -26009, -24134, -19789, -16797, 
    -13758, -8843, -6017, -1372, 5084, 7799, 12712, 16587, 19672, 23062, 
    24526, 27203, 27986, 30752, 30332, 30219, 29454, 29155, 27162, 23895, 
    20311, 18013, 13562, 10034, 7007, -106, -4537, -8276, -10968, -15928, 
    -20954, -22410, -24443, -28140, -27542, -30256, -31587, -29387, -30413, 
    -29102, -25928, -23410, -21286, -18014, -13190, -10665, -6730, -1676, 
    3440, 7090, 11647, 13944, 18984, 22512, 24162, 27977, 28103, 29809, 
    30773, 31113, 29845, 27347, 26898, 24152, 19655, 19029, 13184, 9945, 
    5218, 617, -3946, -8368, -12148, -14490, -18906, -22596, -26183, -26930, 
    -30599, -31066, -30563, -31077, -30928, -29091, -27823, -23911, -20398, 
    -18658, -14643, -9621, -5793, -2089, 4203, 7923, 12320, 14989, 19753, 
    21361, 25086, 28549, 28548, 31366, 29694, 30902, 30107, 28356, 27334, 
    25870, 21364, 17704, 14054, 11496, 7222, 2691, -2627, -7585, -9799, 
    -14490, -17629, -20717, -25514, -26975, -27552, -30080, -30702, -31596, 
    -28456, -29033, -27325, -25639, -21269, -17149, -15304, -10974, -7047, 
    -3149, 1780, 8111, 10414, 15917, 19110, 21551, 24176, 27031, 29141, 
    29425, 31180, 31402, 29286, 28036, 26843, 25155, 22706, 18134, 13900, 
    11722, 7971, 2000, -3801, -6671, -9385, -13112, -19135, -21292, -25935, 
    -26214, -28251, -31394, -30666, -31029, -29801, -29842, -26570, -25891, 
    -22101, -17709, -14987, -11579, -7680, -2841, 1061, 7422, 10446, 13656, 
    17853, 21985, 24923, 25778, 29935, 30841, 31592, 30014, 28601, 29119, 
    28458, 25957, 22610, 19011, 15323, 11723, 6981, 3476, -2172, -6570, 
    -9394, -15629, -17680, -20191, -25923, -24988, -28243, -29848, -30430, 
    -30543, -31109, -28910, -28035, -24152, -22376, -19470, -15334, -12079, 
    -6891, -2685, 1201, 5592, 9796, 13834, 18315, 20899, 23925, 26230, 29604, 
    29037, 29851, 30629, 30304, 29034, 27297, 26191, 22972, 19415, 15677, 
    11041, 8173, 4044, -1361, -5793, -10720, -13110, -18626, -20944, -23954, 
    -24640, -29090, -28820, -31921, -30490, -29955, -29623, -26950, -25547, 
    -22757, -19683, -15604, -12097, -7282, -2706, 320, 5673, 9484, 14941, 
    15958, 19725, 24066, 27172, 29156, 29713, 29442, 30700, 30216, 30552, 
    26684, 24728, 21671, 20230, 15890, 11256, 7553, 4233, -697, -4109, -9083, 
    -13079, -16990, -20463, -24024, -26571, -28106, -31275, -32402, -30947, 
    -30113, -29991, -27493, -25340, -21635, -19340, -16728, -11721, -8936, 
    -4628, -286, 3298, 8890, 13398, 17655, 20589, 23906, 26393, 27397, 29429, 
    30255, 31162, 29227, 28616, 28508, 25962, 22615, 19231, 17138, 11321, 
    7626, 5701, -7, -4777, -9252, -14287, -17290, -20500, -24145, -25984, 
    -27982, -29365, -29966, -30771, -29347, -29258, -28373, -25006, -21839, 
    -19596, -18075, -13509, -7897, -3897, -206, 4622, 7783, 11991, 16744, 
    21426, 24084, 25728, 27558, 30607, 29613, 30305, 30706, 29730, 28932, 
    26418, 23907, 19313, 17034, 12130, 7987, 6341, 948, -3667, -8726, -11130, 
    -16947, -20166, -22829, -25527, -27491, -29502, -31486, -31069, -29037, 
    -29147, -28343, -25486, -22304, -20576, -16652, -13308, -8720, -5532, 
    -568, 4889, 7848, 12322, 16200, 20302, 21543, 25931, 27908, 30810, 28668, 
    30783, 29632, 30058, 27189, 28052, 24970, 20654, 16990, 12832, 9059, 
    6546, 610, -4107, -7103, -12166, -15443, -20590, -24125, -26107, -28211, 
    -29314, -29950, -29398, -30713, -29790, -28324, -26736, -23835, -20708, 
    -18436, -12908, -8362, -5448, -1285, 3452, 7903, 12552, 16294, 19253, 
    22745, 24911, 27414, 30947, 30542, 30568, 30412, 29940, 28117, 25822, 
    23462, 22139, 17440, 14441, 9478, 5269, 1038, -3101, -8213, -12461, 
    -16181, -18402, -23684, -25961, -28125, -30090, -30849, -30010, -31117, 
    -30016, -28154, -25835, -25614, -20405, -19114, -13802, -9714, -5329, 
    -740, 4700, 6414, 10526, 15421, 19871, 21384, 25226, 27026, 29401, 30189, 
    30936, 31169, 30463, 28617, 27804, 25319, 20335, 16453, 15149, 8855, 
    5334, 3121, -3261, -7158, -11122, -15253, -19143, -22532, -26062, -27388, 
    -28322, -30502, -31279, -29414, -30056, -27739, -27232, -24167, -22363, 
    -18342, -15258, -10348, -4664, -1780, 2944, 7389, 10295, 16235, 18395, 
    22274, 25533, 26599, 29273, 30997, 30333, 30849, 31458, 28901, 26248, 
    25140, 21602, 19526, 14920, 11970, 6578, 3266, -1941, -6993, -9894, 
    -13971, -18127, -21902, -24308, -28730, -29104, -29806, -31081, -31008, 
    -28933, -30612, -26272, -26397, -20660, -16984, -14873, -11183, -6845, 
    -2652, 1815, 6370, 10629, 13831, 17815, 21990, 23221, 27150, 27641, 
    29798, 31389, 30048, 29027, 27720, 26418, 24981, 20660, 17802, 13731, 
    11127, 6304, 1234, -2193, -6757, -10280, -14442, -18686, -22411, -23849, 
    -26692, -26996, -29076, -30732, -30449, -30082, -28561, -26248, -24243, 
    -23401, -18758, -15413, -12042, -6360, -2041, 2075, 7025, 10581, 14516, 
    18111, 22061, 24310, 26821, 27671, 28610, 31870, 29365, 30084, 28740, 
    28358, 25436, 23379, 20205, 15176, 12695, 6994, 1689, -920, -5520, 
    -11169, -13640, -17909, -21820, -24382, -26495, -30115, -29169, -31632, 
    -29838, -29984, -29482, -26780, -24255, -21435, -18718, -14651, -11572, 
    -7531, -2614, 580, 6170, 10649, 13305, 17656, 20301, 23742, 26033, 26900, 
    30336, 30719, 31193, 29460, 28977, 27546, 24018, 22454, 19026, 15968, 
    10719, 8013, 3569, -823, -4980, -8866, -13555, -18078, -21014, -23643, 
    -26483, -28353, -31178, -30440, -30472, -30600, -29369, -26301, -25148, 
    -23608, -19476, -15134, -11545, -6832, -3434, 459, 5493, 9565, 13660, 
    18044, 21094, 22099, 26365, 28372, 30090, 29699, 31283, 29300, 30030, 
    28714, 26647, 23090, 19144, 16353, 12491, 8478, 4548, 479, -4772, -9303, 
    -12353, -17264, -20772, -23297, -26294, -28170, -28814, -30318, -30838, 
    -30913, -29491, -28896, -26973, -22572, -20664, -16946, -11922, -6770, 
    -2552, -603, 5328, 10335, 13737, 16741, 19910, 24327, 26975, 27960, 
    29377, 30683, 31221, 30756, 29423, 28057, 27561, 21594, 20135, 16401, 
    11185, 9643, 4983, -515, -4096, -7661, -13544, -15911, -19027, -23634, 
    -25825, -29555, -30449, -31235, -30906, -30620, -30725, -28317, -25206, 
    -23238, -20568, -16764, -12223, -8905, -5907, 767, 3746, 10223, 11542, 
    16768, 20394, 22458, 26382, 26462, 30322, 30507, 30963, 31025, 28934, 
    28020, 25678, 22326, 21196, 17678, 12404, 9015, 3636, 597, -3827, -7377, 
    -12296, -16169, -20256, -24583, -24660, -26799, -31091, -30514, -31083, 
    -30414, -30314, -27459, -24759, -25099, -20177, -17165, -13422, -7316, 
    -3706, -991, 4901, 7754, 13530, 16451, 19866, 24467, 25704, 27617, 29439, 
    30876, 30612, 29625, 28848, 28249, 26851, 23079, 21714, 16630, 13609, 
    9553, 6483, 306, -5211, -8515, -11391, -15856, -20098, -23333, -25887, 
    -27252, -29560, -29676, -31645, -30827, -30795, -29181, -25332, -24458, 
    -21899, -16919, -14440, -7854, -5557, -502, 3548, 7290, 11583, 16165, 
    19600, 22407, 25563, 27858, 30345, 30313, 29767, 30282, 29478, 29683, 
    26210, 23303, 21338, 16936, 14164, 8917, 5902, 1943, -3248, -6375, 
    -10467, -14580, -17678, -22149, -24844, -27802, -28661, -30104, -30724, 
    -31534, -29955, -27603, -26684, -24919, -20969, -17377, -15006, -8984, 
    -4198, -2866, 2138, 7556, 12013, 14906, 19065, 22233, 24473, 26948, 
    28758, 29211, 30276, 30698, 30280, 28437, 26944, 24042, 21513, 18042, 
    15155, 9644, 6009, 2766, -1918, -8037, -11278, -14516, -18676, -23078, 
    -25565, -28764, -28057, -31164, -30546, -31160, -28764, -29040, -26605, 
    -25046, -22643, -17649, -15079, -10345, -5802, -879, 4075, 7193, 11577, 
    14123, 19411, 22634, 26441, 26482, 28132, 30510, 30719, 29283, 30419, 
    28627, 27503, 25475, 22645, 16805, 14856, 11312, 6710, 1936, -734, -6663, 
    -11799, -15830, -17531, -21184, -24666, -26887, -29295, -30716, -30553, 
    -29518, -30099, -28736, -27163, -25932, -22906, -19990, -14783, -12057, 
    -6316, -1310, 2632, 5914, 11885, 15237, 18672, 22513, 24767, 25950, 
    27586, 30185, 30125, 31456, 28824, 29452, 25804, 25890, 20769, 18399, 
    15370, 11966, 6683, 4109, -3173, -6813, -10507, -14548, -17024, -21603, 
    -24884, -26327, -27712, -30031, -30729, -30318, -30160, -28872, -27828, 
    -25668, -20800, -18193, -14818, -10640, -7191, -3087, 455, 5200, 10009, 
    14751, 18178, 20206, 24228, 26105, 28777, 30565, 31220, 30139, 29631, 
    29273, 28783, 24068, 23176, 19490, 15167, 10973, 7829, 3119, -329, -5537, 
    -11181, -14488, -19239, -22104, -23812, -26787, -30102, -29458, -29582, 
    -30770, -29807, -27935, -26844, -25939, -23450, -19494, -15403, -12904, 
    -8252, -3169, 1377, 4605, 9973, 14396, 18720, 20010, 23904, 25988, 28693, 
    29823, 29552, 30503, 29616, 29225, 28413, 25070, 22743, 20102, 16687, 
    11420, 7577, 2093, -1679, -5051, -10664, -14449, -16956, -21387, -24524, 
    -27698, -28149, -30418, -30375, -31103, -28899, -29986, -28936, -25514, 
    -22423, -18378, -17663, -11471, -8847, -4849, -192, 5350, 10435, 15257, 
    16279, 20713, 22842, 25314, 27502, 30454, 29364, 29515, 30417, 28536, 
    25838, 24160, 22290, 19445, 15987, 12284, 8191, 3934, -284, -6470, 
    -10465, -13351, -16680, -22039, -23340, -25103, -28726, -30101, -30381, 
    -30974, -30838, -29173, -26285, -25877, -23032, -19466, -17724, -11278, 
    -9459, -3238, -1213, 5674, 9384, 13366, 16656, 19180, 23291, 26379, 
    28133, 29746, 31781, 31927, 30838, 29116, 27801, 25218, 23494, 20962, 
    15183, 13741, 10043, 5192, -633, -4024, -9371, -11975, -17411, -20388, 
    -23370, -26523, -28302, -30254, -30012, -30227, -30101, -29673, -26628, 
    -27633, -23642, -20067, -16839, -13851, -7994, -4234, 344, 3447, 8346, 
    12268, 16607, 19320, 23735, 25742, 27626, 29206, 30250, 30789, 30327, 
    29909, 27048, 25638, 23069, 19415, 16958, 12252, 8278, 5025, 1584, -5019, 
    -8258, -11315, -17132, -20146, -23248, -25495, -28668, -28977, -30823, 
    -30168, -29408, -31183, -27428, -25447, -22601, -20425, -18400, -11758, 
    -10150, -3218, -748, 4152, 8327, 13767, 15591, 19145, 23090, 24884, 
    27384, 29906, 30784, 32190, 30025, 30504, 28875, 25990, 22078, 20511, 
    16608, 14608, 8458, 5864, 379, -3650, -7560, -11407, -15902, -19339, 
    -23872, -27121, -27870, -28533, -30079, -29476, -30181, -28467, -27472, 
    -26795, -23784, -20853, -17645, -14643, -9175, -4995, -373, 3090, 7220, 
    12027, 15337, 18754, 24434, 24800, 29392, 29273, 30915, 30915, 31375, 
    30353, 28611, 25614, 23092, 21188, 16948, 12633, 8643, 3907, 645, -3878, 
    -7216, -10650, -15520, -19095, -21999, -23578, -27165, -30053, -31370, 
    -30316, -29301, -30847, -27264, -26510, -23139, -21286, -17151, -13566, 
    -8876, -5392, -50, 4068, 8375, 10551, 15084, 20030, 20742, 24026, 26066, 
    29066, 29232, 30323, 30384, 31395, 29445, 27422, 24924, 20490, 17450, 
    13730, 10169, 4369, 39, -1995, -7061, -11427, -15818, -19313, -21838, 
    -24542, -26834, -28722, -30447, -31347, -29969, -29684, -27995, -26495, 
    -24889, -21338, -17511, -15787, -12118, -6361, -1046, 2557, 7332, 11441, 
    16011, 18112, 22909, 25870, 26575, 29244, 30558, 30639, 30796, 30492, 
    28629, 26688, 24641, 22204, 18442, 14611, 10421, 7105, 1438, -2689, 
    -7726, -10689, -13365, -18728, -21857, -23935, -28279, -28890, -30696, 
    -30920, -29723, -30499, -29022, -26780, -25185, -20823, -18234, -15897, 
    -11761, -6309, -879, 1463, 5235, 10000, 15500, 19549, 21189, 23801, 
    28251, 27213, 29273, 30364, 31558, 28841, 28511, 28481, 24939, 21447, 
    19012, 15332, 10698, 7301, 1595, -2579, -6204, -10438, -14268, -17354, 
    -21499, -23544, -26913, -28561, -29937, -30777, -30327, -31148, -27804, 
    -26799, -25386, -20772, -19132, -14094, -11240, -6454, -2003, 1115, 6251, 
    12187, 14484, 19192, 20016, 23253, 28330, 28213, 29059, 29150, 31253, 
    29274, 29543, 27716, 23520, 21872, 18289, 15373, 11908, 5375, 2639, 
    -1430, -7416, -11225, -14415, -17536, -20629, -24079, -26888, -29650, 
    -29095, -30496, -30649, -31593, -30017, -27105, -26399, -23002, -20233, 
    -15493, -12572, -6020, -1513, 2366, 6713, 10758, 14620, 17384, 21800, 
    24101, 25473, 28018, 29134, 30179, 32065, 31095, 28672, 27556, 25318, 
    21285, 20136, 16982, 11725, 6703, 3646, -2208, -5194, -9993, -13252, 
    -17644, -21405, -24483, -27191, -29284, -29707, -32161, -29733, -28594, 
    -29084, -27750, -25445, -22384, -20263, -16319, -12658, -7622, -2749, 
    1461, 7096, 9520, 14952, 17253, 21911, 24018, 26653, 28216, 29422, 30399, 
    31603, 30289, 28888, 26252, 25090, 22051, 19863, 16390, 12938, 9170, 
    3381, -1881, -6502, -8151, -14435, -16046, -20900, -23689, -25678, 
    -29068, -29939, -29959, -30385, -30337, -28932, -27091, -24969, -22913, 
    -19467, -17817, -11682, -7593, -4031, 1890, 6015, 10161, 13949, 15668, 
    18696, 23270, 26342, 27635, 31373, 29718, 29772, 28938, 28845, 28758, 
    26425, 23512, 21561, 15907, 11855, 9701, 4511, -223, -5604, -8453, 
    -13360, -17428, -21730, -22839, -27520, -27366, -28895, -31364, -31552, 
    -28786, -30306, -26947, -26488, -25134, -21003, -17288, -12324, -10125, 
    -5387, 489, 3470, 8319, 12954, 17049, 19165, 23238, 26009, 28880, 30484, 
    29977, 31280, 30579, 29511, 28722, 27262, 23649, 19945, 16111, 11496, 
    10269, 5663, 634, -3425, -8500, -12393, -16350, -19822, -24121, -26890, 
    -27610, -29463, -30210, -30925, -30816, -29236, -26568, -24943, -23750, 
    -21151, -17141, -11673, -8844, -4112, 276, 3587, 8600, 11433, 17528, 
    18886, 22463, 25953, 28796, 27818, 31507, 30165, 31156, 28644, 28821, 
    26273, 24131, 20597, 17250, 12932, 9846, 4656, 48, -4067, -8293, -11323, 
    -16225, -19892, -22319, -24149, -27646, -29959, -30792, -31906, -29603, 
    -29602, -26815, -26818, -23219, -19427, -16907, -13034, -9702, -6346, 
    -523, 3275, 8014, 11395, 15832, 20290, 21960, 26334, 27912, 29339, 31145, 
    30765, 30872, 28396, 27619, 26827, 23227, 20859, 18234, 13898, 9452, 
    5138, 2204, -4059, -6657, -9957, -15769, -18357, -22093, -25999, -27069, 
    -29898, -29690, -29685, -30895, -30902, -28986, -27984, -24681, -21434, 
    -17425, -14938, -11579, -6105, -515, 3728, 8070, 11658, 15914, 19383, 
    22249, 25803, 27706, 29221, 31415, 29333, 30033, 28848, 27286, 26855, 
    23781, 21311, 19011, 14703, 8962, 5241, 1506, -1499, -7829, -11204, 
    -15360, -19781, -22729, -24776, -27277, -28461, -31120, -30842, -31204, 
    -28185, -28306, -26962, -23084, -22753, -17729, -14215, -10702, -5615, 
    -1244, 1985, 6969, 11320, 15486, 19186, 21858, 23513, 27418, 27664, 
    31731, 30140, 30199, 28798, 27239, 27689, 25144, 23193, 18585, 15866, 
    11173, 7133, 2451, -1816, -7185, -11032, -16108, -16888, -20858, -24834, 
    -26167, -29264, -29737, -30675, -29507, -29942, -27328, -27048, -24242, 
    -22458, -18239, -15397, -9440, -6977, -2144, 1466, 6828, 10799, 15453, 
    17411, 23103, 24553, 28117, 28786, 30796, 31956, 30997, 29968, 28949, 
    28779, 26287, 21418, 18364, 15293, 11816, 8598, 2084, -685, -6575, 
    -10300, -13586, -17678, -21423, -24752, -26924, -30091, -28882, -31839, 
    -29722, -29858, -28457, -27242, -25438, -21597, -18640, -15334, -11978, 
    -8199, -3743, 2564, 6848, 10461, 13304, 18941, 21840, 23483, 26603, 
    30251, 30430, 31517, 30298, 29074, 28618, 27774, 26489, 22397, 19208, 
    16597, 10431, 7712, 1141, -470, -4909, -11532, -15372, -18643, -21946, 
    -25261, -27864, -28648, -30205, -30415, -30064, -29567, -30830, -29218, 
    -25683, -24085, -18153, -15511, -12691, -7502, -1630, 2482, 5692, 10692, 
    15459, 16705, 21995, 24351, 26275, 27956, 31157, 30411, 31725, 30768, 
    28784, 27886, 23586, 22484, 19916, 15584, 11054, 7063, 3019, 53, -6691, 
    -10322, -14365, -17308, -20586, -24080, -26372, -28793, -31509, -31621, 
    -30373, -30805, -29629, -27287, -24778, -22530, -20208, -15410, -12241, 
    -6148, -2292, 410, 5329, 9546, 14135, 16780, 20464, 23267, 26162, 28014, 
    29239, 29801, 30251, 30954, 30022, 29218, 25350, 22872, 21075, 15379, 
    12695, 7750, 2564, -61, -3858, -8633, -13129, -17523, -20793, -24815, 
    -25252, -29787, -28985, -29103, -30236, -29990, -29507, -28006, -24823, 
    -23430, -20091, -18026, -12744, -7888, -2525, 272, 4665, 9620, 14290, 
    18298, 20662, 23542, 26952, 29098, 30736, 30510, 32343, 30707, 29924, 
    29327, 25377, 22631, 20638, 15817, 12942, 8727, 3510, -441, -4727, -7181, 
    -13732, -17699, -20922, -24990, -25987, -27657, -29652, -29374, -31431, 
    -28829, -29305, -27498, -24437, -22316, -20303, -16417, -11513, -9164, 
    -4267, 1329, 4366, 8901, 11433, 16199, 20329, 23135, 24865, 27614, 30061, 
    30666, 30870, 30289, 29375, 29133, 27119, 22905, 20686, 15950, 13011, 
    9550, 4345, -310, -5132, -8046, -11959, -15125, -19855, -22036, -24399, 
    -28744, -29292, -30138, -31199, -29883, -30615, -28143, -27057, -24081, 
    -19178, -17703, -12766, -9229, -4720, -44, 3406, 8616, 11787, 17106, 
    20249, 22984, 24495, 28226, 28894, 28684, 30093, 32363, 30555, 26679, 
    26565, 24806, 20085, 18008, 14541, 10705, 5077, 156, -2801, -8011, 
    -13400, -16575, -19234, -21727, -26247, -26780, -29735, -30156, -31505, 
    -30641, -31255, -28549, -26401, -24929, -21387, -16966, -14536, -9120, 
    -4384, 641, 2901, 6990, 11063, 15810, 18832, 23197, 25878, 28627, 29345, 
    31615, 31285, 31156, 30582, 27885, 25565, 24874, 22222, 17275, 13974, 
    9543, 5718, 1824, -2509, -7991, -11140, -14419, -18410, -23764, -24428, 
    -27095, -29452, -31853, -31317, -29779, -30922, -29536, -27424, -23955, 
    -21692, -18334, -15543, -11078, -5899, -681, 1711, 6126, 9754, 16027, 
    19862, 20700, 26637, 27150, 28542, 31889, 31462, 30259, 28267, 29636, 
    27171, 23657, 20862, 16735, 13909, 11297, 4297, 379, -2272, -7344, 
    -12521, -15711, -19582, -21458, -25281, -26648, -30136, -28851, -31011, 
    -31931, -29512, -28972, -26915, -23567, -20315, -17645, -14732, -10699, 
    -5591, -785, 3175, 6736, 10406, 15632, 18364, 21944, 25584, 25986, 28316, 
    30232, 31372, 30795, 30393, 29559, 26605, 24079, 20523, 17919, 14567, 
    10442, 6053, 965, -3355, -6482, -10049, -13435, -17892, -21331, -24803, 
    -27532, -30204, -28975, -31470, -31585, -31804, -28732, -27633, -24530, 
    -21259, -18648, -15214, -9015, -4931, -2908, 3900, 6272, 10515, 12819, 
    17054, 22088, 25827, 26178, 28838, 30885, 31302, 30782, 30275, 29511, 
    27000, 25454, 21351, 19043, 14468, 10459, 6868, 3204, -3272, -6067, 
    -9120, -14617, -17257, -20450, -24250, -27681, -28480, -31083, -31671, 
    -30497, -31207, -28551, -25727, -25430, -23388, -18597, -15087, -11441, 
    -6934, -1874, 1497, 6288, 10516, 13708, 19038, 22568, 23795, 25989, 
    27600, 30502, 30312, 29806, 30567, 28846, 27452, 24767, 21029, 18471, 
    16462, 10058, 7304, 3225, -926, -6676, -9617, -14490, -19481, -21166, 
    -22899, -25636, -28375, -29629, -30703, -30325, -30964, -30085, -27780, 
    -24527, -21675, -19594, -16216, -11659, -7224, -2698, 1806, 5720, 9599, 
    14193, 18021, 20966, 24985, 26560, 29575, 29885, 30806, 31298, 30575, 
    28874, 28073, 25255, 22018, 19672, 15776, 12241, 8677, 2953, -313, -5106, 
    -9343, -11978, -17738, -21083, -22945, -25832, -28937, -29386, -30211, 
    -29639, -30815, -29778, -27539, -25989, -22559, -19034, -16023, -12936, 
    -6949, -4741, 401, 5332, 10768, 14358, 17228, 21783, 22289, 25435, 27733, 
    29690, 30947, 30692, 30582, 29034, 26790, 25075, 22763, 20092, 14795, 
    11510, 6699, 3396, -1078, -4718, -9906, -13987, -15820, -20992, -23237, 
    -26848, -28059, -29592, -31557, -31136, -29725, -29730, -27822, -25255, 
    -22842, -19978, -15314, -11025, -6750, -3821, 518, 3900, 9857, 12968, 
    16714, 19500, 24381, 25133, 27778, 29535, 30216, 30340, 29867, 30383, 
    29262, 26828, 22020, 20977, 17903, 13610, 7941, 3259, 693, -4939, -9473, 
    -12970, -16757, -19701, -23203, -25715, -28113, -29939, -29524, -31842, 
    -29097, -29598, -27928, -25956, -24085, -18686, -16845, -12562, -9004, 
    -4506, -594, 3637, 9343, 13121, 17702, 21979, 23350, 25693, 27693, 30493, 
    30558, 32523, 31998, 30810, 29156, 27226, 22701, 21110, 16142, 13995, 
    8906, 4847, -428, -4814, -7674, -13589, -17759, -20998, -23387, -24634, 
    -28463, -29290, -31814, -31301, -30609, -28704, -27087, -26242, -22196, 
    -19853, -16655, -13131, -8870, -5727, 1389, 3476, 8328, 11893, 16704, 
    18962, 24062, 26462, 27899, 29350, 29312, 30061, 30211, 29489, 26803, 
    27583, 23569, 21757, 16076, 14654, 9581, 3949, 412, -5116, -7106, -13194, 
    -15372, -19733, -22583, -24582, -26244, -28756, -30418, -32469, -30688, 
    -28633, -28391, -26949, -22786, -19270, -19141, -12719, -11103, -6279, 
    -621, 3494, 7604, 12786, 14695, 18095, 22484, 25426, 29269, 27910, 31058, 
    31411, 29230, 30826, 27940, 26374, 24043, 21395, 17630, 15211, 9019, 
    6421, 563, -5124, -7549, -11962, -16927, -19470, -23211, -25244, -27324, 
    -29435, -31786, -31428, -31001, -30497, -27670, -24743, -23960, -21985, 
    -17690, -12256, -10419, -4984, -1379, 3072, 8389, 12457, 16116, 20224, 
    22404, 25854, 28706, 28206, 29840, 30862, 29678, 30470, 28364, 26836, 
    22707, 21616, 18670, 15178, 10157, 5429, 761, -1811, -8441, -11829, 
    -15585, -19539, -21662, -25421, -26694, -28693, -29180, -30921, -31935, 
    -30709, -28103, -27091, -22931, -22055, -18523, -14501, -11225, -5246, 
    -842, 2408, 6696, 10269, 13750, 17540, 22509, 24954, 25900, 29179, 29769, 
    30718, 31418, 29941, 27240, 26608, 25028, 20894, 17136, 13794, 10534, 
    6798, 1929, -3128, -6001, -10121, -16352, -18129, -22423, -23919, -28173, 
    -28586, -29934, -29109, -30461, -28935, -28124, -26922, -25046, -21652, 
    -18393, -15709, -10889, -6456, -803, 1635, 6643, 9562, 13950, 18413, 
    20471, 25371, 27654, 28697, 30165, 29956, 30615, 31376, 28277, 26297, 
    23396, 21459, 18533, 15195, 10022, 7211, 3424, -966, -6408, -11117, 
    -14036, -19714, -21604, -24825, -25765, -29237, -30706, -30168, -30139, 
    -30694, -29245, -26367, -24151, -21535, -17751, -15278, -12675, -7569, 
    -3980, 1374, 6082, 10710, 12786, 19311, 20432, 22865, 28412, 28980, 
    29629, 29886, 31813, 29823, 30691, 27861, 25255, 22080, 19605, 15625, 
    12233, 6928, 2754, -956, -6400, -10932, -14420, -17764, -22051, -25771, 
    -26274, -28502, -30170, -30131, -32170, -29052, -28802, -25982, -24280, 
    -21689, -18838, -16145, -11929, -7269, -1901, 870, 5049, 9480, 14455, 
    16998, 22510, 22670, 25261, 27923, 29652, 31562, 30414, 30336, 29401, 
    28607, 24395, 22035, 18738, 15407, 11854, 6457, 4523, -293, -5467, 
    -10060, -13170, -18691, -19779, -22222, -25806, -27977, -30510, -30416, 
    -30831, -29573, -28756, -28081, -26788, -22462, -20405, -15981, -13873, 
    -8513, -2167, 1468, 5977, 8527, 12294, 18353, 21543, 22322, 26642, 29374, 
    29948, 28800, 29634, 29564, 28348, 28319, 24225, 22640, 20043, 16836, 
    12558, 8573, 3612, -1016, -4926, -10873, -14110, -17746, -20059, -23931, 
    -25597, -27820, -29696, -30467, -30773, -31054, -29421, -26941, -25816, 
    -22307, -20656, -16335, -12981, -7997, -3719, -108, 3662, 8974, 14002, 
    16616, 20888, 23144, 25581, 27674, 29144, 29897, 31709, 31881, 30000, 
    28110, 25578, 22469, 19466, 15749, 11434, 8194, 2878, -463, -3602, -7824, 
    -12983, -16168, -20943, -25213, -26959, -27882, -29791, -30581, -31750, 
    -32007, -29507, -26706, -25563, -23783, -18756, -16728, -11754, -9454, 
    -5614, -1488, 5893, 9268, 11942, 15770, 18529, 21832, 24904, 26669, 
    30794, 32171, 30566, 30023, 30208, 26863, 25707, 23748, 19555, 15941, 
    13981, 8966, 5090, 308, -3690, -9244, -12799, -15540, -20590, -22369, 
    -24760, -27397, -30192, -31358, -31349, -29848, -28592, -28672, -26982, 
    -22539, -20713, -17021, -12733, -8270, -6613, -398, 4974, 7443, 11296, 
    15557, 19901, 22912, 25047, 27157, 29501, 29102, 31210, 29938, 30062, 
    28831, 26482, 22706, 20437, 17818, 11729, 10239, 4375, 1215, -3523, 
    -7132, -10524, -14544, -19268, -21875, -26672, -29040, -29126, -31674, 
    -32071, -30310, -30087, -28782, -24660, -24003, -20471, -18286, -12959, 
    -9621, -5195, -911, 3179, 8729, 12993, 15424, 19152, 21570, 24986, 29403, 
    29577, 30572, 29752, 30456, 29774, 27438, 26582, 22776, 20000, 18227, 
    13770, 9065, 6343, 1516, -2470, -7695, -11472, -15936, -19871, -21826, 
    -24294, -27896, -29541, -29098, -31421, -30098, -31085, -27278, -27515, 
    -23636, -20355, -16435, -14471, -8247, -5940, -725, 2762, 7403, 11741, 
    16082, 20705, 22917, 24607, 27365, 28217, 30128, 29895, 29691, 29842, 
    27468, 26787, 23983, 21389, 17587, 13670, 9525, 6904, 1580, -2442, -6007, 
    -11094, -16504, -19223, -21106, -25037, -28177, -27966, -30499, -31913, 
    -31166, -30164, -29100, -25561, -24581, -20929, -17688, -13895, -11439, 
    -6938, -2276, 1278, 7040, 12973, 14697, 19541, 23854, 24681, 25794, 
    29325, 30096, 29758, 30927, 29799, 29821, 27021, 25439, 20576, 18738, 
    14204, 12099, 7526, 2261, -4057, -7792, -12315, -15016, -19316, -21250, 
    -26164, -27334, -29135, -30106, -30185, -32126, -29878, -29237, -27123, 
    -24710, -21023, -17589, -15864, -12011, -5171, -2932, 1997, 5265, 10448, 
    13248, 17919, 21637, 26322, 25723, 29602, 29263, 31559, 30573, 30342, 
    29427, 26795, 25436, 22576, 19494, 14680, 12298, 6685, 1785, -1326, 
    -7005, -10238, -14810, -17605, -21022, -24315, -25950, -28054, -30820, 
    -31862, -31822, -29987, -27715, -26572, -25548, -22164, -17473, -15808, 
    -10325, -6287, -1252, 495, 7208, 10031, 12757, 18280, 21978, 24129, 
    26978, 27498, 29506, 31359, 30851, 31115, 28163, 27102, 24904, 22218, 
    20251, 15270, 10448, 8326, 3869, -2114, -6643, -10443, -13276, -19235, 
    -21206, -25513, -26445, -29487, -29056, -29981, -31441, -30916, -29520, 
    -28900, -24173, -23763, -19999, -16269, -11537, -7632, -3690, -94, 5410, 
    10196, 12887, 17609, 21390, 24139, 28249, 27784, 30292, 31649, 30649, 
    29922, 29867, 27937, 24585, 23294, 19437, 16951, 11282, 6509, 3928, -497, 
    -5071, -10778, -13192, -18595, -22091, -24558, -26449, -29044, -29269, 
    -30536, -31269, -29901, -29456, -28156, -25041, -22670, -19372, -14571, 
    -11691, -8989, -2663, 434, 3945, 9272, 12984, 18826, 20131, 24331, 26682, 
    30083, 30444, 30127, 29485, 29241, 28967, 27289, 25594, 22233, 18217, 
    15160, 13332, 6505, 2040, -116, -4191, -10911, -13186, -16390, -21452, 
    -23777, -26242, -27811, -29765, -29954, -31841, -31253, -30543, -27162, 
    -25097, -22935, -19224, -16222, -13415, -8247, -3699, 1988, 3198, 10265, 
    12650, 18328, 19123, 23813, 26707, 26637, 29436, 31328, 30981, 30601, 
    29754, 27406, 25594, 24328, 18860, 18198, 13376, 8469, 3747, 826, -4535, 
    -8704, -14208, -15787, -20801, -23119, -27000, -28016, -28469, -29934, 
    -29736, -29870, -29840, -28573, -26569, -22737, -19926, -17702, -12977, 
    -7282, -4443, 478, 3580, 7680, 13744, 16407, 20275, 23761, 25037, 28753, 
    30139, 30523, 30307, 30398, 28247, 26977, 26184, 24510, 20685, 18525, 
    12335, 10061, 4823, 786, -4670, -8788, -10948, -15173, -18501, -22367, 
    -27535, -27247, -29166, -29488, -31337, -30233, -30030, -28358, -24999, 
    -23182, -19956, -16975, -13092, -8596, -3350, -800, 2941, 6923, 12220, 
    15495, 18540, 22010, 26309, 28598, 29423, 32156, 32230, 30784, 30488, 
    28374, 26149, 24536, 21358, 17978, 12930, 10547, 4720, 1146, -3090, 
    -8249, -10969, -16955, -20861, -21944, -25457, -28707, -28781, -31059, 
    -30177, -28975, -30122, -27271, -26885, -23967, -19724, -16664, -12872, 
    -10509, -6877, -1668, 3182, 8212, 12756, 15988, 18752, 22741, 27111, 
    28568, 29665, 30836, 29821, 30631, 29522, 28861, 27869, 24456, 19632, 
    17524, 12955, 8546, 5901, 2273, -2504, -8109, -11539, -15452, -18745, 
    -22191, -26553, -26667, -28487, -29630, -31385, -30940, -30229, -27248, 
    -27028, -23429, -21960, -18050, -13834, -8658, -6100, -486, 2833, 7509, 
    11844, 15482, 18936, 22339, 26760, 27383, 28350, 30735, 29305, 31566, 
    28576, 26866, 25722, 25231, 19556, 16242, 13611, 10995, 6886, 3000, 
    -2956, -7785, -11945, -14436, -19075, -21261, -25536, -25476, -29742, 
    -29540, -29992, -28837, -29056, -28295, -27150, -24906, -20973, -17463, 
    -14717, -11593, -6271, -1728, 2688, 6684, 9517, 15270, 18416, 21981, 
    25911, 27085, 30556, 29500, 31669, 29895, 30673, 29709, 27061, 25040, 
    22540, 17587, 15685, 10484, 6445, 1542, -1272, -7789, -10747, -14049, 
    -18525, -21213, -24179, -26002, -30808, -30680, -30550, -29998, -29667, 
    -29747, -27808, -26095, -21506, -18711, -14568, -10210, -8279, -726, 
    1279, 5673, 10886, 14725, 19568, 22242, 24694, 27899, 27896, 30853, 
    29347, 29449, 29722, 27803, 26050, 24833, 22804, 19640, 15275, 10752, 
    7328, 1772, -2633, -5180, -11293, -15722, -18493, -21027, -24682, -28094, 
    -29595, -30717, -32205, -31169, -30165, -30078, -26619, -26382, -23121, 
    -18805, -16308, -11815, -6145, -1943, 1514, 5858, 11635, 14888, 19419, 
    23060, 24246, 26487, 29438, 29469, 29613, 30595, 30276, 28619, 27547, 
    25603, 21798, 18449, 16478, 10818, 7833, 1519, -1553, -6957, -8281, 
    -13947, -17265, -19805, -23524, -27722, -28928, -29760, -29874, -30691, 
    -30429, -29117, -26676, -24952, -22556, -19408, -15235, -10515, -8319, 
    -2727, 1263, 5150, 10248, 13814, 16254, 21246, 23871, 27310, 28016, 
    30373, 30843, 30436, 29871, 27982, 27745, 25185, 22679, 18691, 14470, 
    10061, 8438, 3687, -282, -7029, -9784, -13825, -18190, -22397, -23288, 
    -26257, -28690, -29685, -29432, -31468, -29602, -28839, -27983, -25194, 
    -22382, -19368, -15229, -10609, -7010, -4785, 983, 4267, 8086, 13074, 
    15798, 21141, 23549, 26319, 28247, 30918, 29402, 32244, 31977, 29449, 
    27368, 26238, 22384, 20482, 16961, 10828, 6300, 5528, -443, -4481, -9241, 
    -12156, -16978, -20262, -23604, -26618, -28193, -30038, -30432, -30808, 
    -29901, -30732, -27129, -26016, -22677, -19356, -16292, -13491, -8216, 
    -2814, -833, 4734, 8974, 12144, 17412, 21450, 22063, 25231, 29355, 29486, 
    31865, 31074, 29306, 30183, 28827, 26214, 22624, 19361, 14627, 12825, 
    8684, 4908, -1037, -4834, -10400, -14008, -16674, -19450, -22274, -26042, 
    -28993, -30273, -30605, -30185, -31206, -29771, -27175, -25281, -24836, 
    -21206, -16156, -12855, -7849, -4690, -1017, 4475, 8585, 11972, 17343, 
    21017, 22424, 25899, 28885, 29805, 31768, 30004, 31355, 29641, 29017, 
    26331, 24870, 21284, 15200, 14740, 8984, 4150, 1155, -4304, -8063, 
    -10891, -17884, -20481, -22743, -24868, -26576, -28587, -28969, -31884, 
    -31942, -30244, -28582, -25690, -24205, -19930, -16300, -11737, -9149, 
    -3603, -1129, 2625, 8617, 12294, 17317, 18301, 23198, 24206, 27897, 
    31198, 28633, 30611, 31186, 30033, 27160, 26404, 24829, 20236, 18769, 
    13496, 8921, 5625, 978, -3686, -8153, -11909, -15281, -20094, -22594, 
    -24154, -27765, -29000, -31332, -30303, -30476, -30992, -28420, -27529, 
    -22642, -21499, -16754, -12842, -9492, -5050, 153, 3847, 9081, 12287, 
    15107, 18137, 22957, 24818, 27868, 29994, 30966, 30729, 30037, 28484, 
    28274, 27000, 23953, 20054, 17847, 14641, 9129, 6829, 983, -3304, -7491, 
    -11246, -14054, -19311, -21978, -25719, -27801, -29505, -31014, -30942, 
    -30859, -30553, -29754, -25815, -24055, -22243, -19195, -13256, -9058, 
    -5751, -1384, 4702, 7903, 10789, 16052, 18561, 22298, 24386, 27128, 
    30162, 29596, 29526, 30368, 30116, 28700, 25243, 22943, 20768, 18348, 
    15054, 10942, 4724, 1791, -4272, -7077, -12504, -15751, -18370, -20871, 
    -24915, -28746, -28186, -30898, -31019, -31577, -30845, -28212, -25388, 
    -24631, -21772, -18850, -13220, -12209, -6083, -3039, 866, 7793, 11833, 
    14910, 18545, 23431, 25349, 28475, 30156, 30808, 32052, 30333, 31483, 
    28289, 25728, 24503, 21965, 17306, 14318, 9905, 5408, 1703, -2463, -6418, 
    -10773, -14297, -18002, -20687, -25230, -27245, -29821, -29007, -31658, 
    -30342, -29690, -28188, -27363, -24884, -22771, -18265, -13761, -9928, 
    -7456, -2645, 1681, 7097, 10256, 16086, 19413, 21516, 25934, 26846, 
    28699, 28708, 30022, 31396, 28780, 28565, 27575, 25883, 21770, 18987, 
    15885, 10186, 8031, 3553, -2408, -6140, -10169, -15856, -17278, -20567, 
    -24256, -28064, -27705, -29853, -31136, -29355, -29352, -28426, -27713, 
    -26678, -21581, -18245, -14789, -11323, -8223, -2623, 1439, 7640, 11844, 
    14528, 17989, 22701, 23247, 27629, 28133, 29607, 30665, 29902, 31408, 
    28406, 26591, 26489, 23108, 19421, 16112, 11286, 7672, 3635, -562, -5229, 
    -10763, -12509, -17788, -21919, -25390, -25061, -28726, -30985, -30275, 
    -31338, -30031, -27539, -28001, -24891, -20631, -18985, -15623, -11478, 
    -7865, -2857, 704, 4604, 10182, 13044, 18685, 20894, 23697, 27540, 29523, 
    29244, 30689, 31485, 30349, 28994, 26619, 25279, 22012, 19593, 16099, 
    11766, 7429, 3416, -191, -6543, -9593, -12796, -18585, -21780, -22816, 
    -25407, -28376, -29498, -30532, -30234, -31606, -28057, -27174, -24820, 
    -21924, -19762, -16017, -12277, -7756, -1836, 1906, 5063, 9700, 11937, 
    17938, 22615, 23746, 28056, 29201, 30370, 30566, 30007, 32118, 28537, 
    27124, 25469, 22630, 20653, 17534, 12476, 8668, 3309, -1447, -3378, 
    -9942, -12472, -15502, -20269, -23911, -25693, -29034, -28982, -30665, 
    -29593, -31983, -29311, -27434, -25111, -22946, -21033, -15722, -12607, 
    -8540, -4119, 548, 5227, 9344, 13695, 17255, 18872, 23231, 26996, 26503, 
    30668, 30856, 30722, 32005, 28185, 27752, 27058, 22602, 18664, 16071, 
    13474, 6601, 3713, 291, -5387, -7780, -14377, -16504, -20759, -23522, 
    -25474, -27597, -29486, -31613, -30348, -29812, -28571, -26998, -26420, 
    -22799, -21215, -16453, -12656, -7989, -4933, -756, 4119, 9107, 13584, 
    16372, 20735, 22641, 25145, 29061, 29631, 29953, 32119, 31526, 29657, 
    28531, 26680, 23222, 20212, 17572, 14347, 10641, 5582, 29, -2787, -7851, 
    -13754, -16703, -18866, -21521, -25725, -28916, -29646, -30245, -30738, 
    -29623, -28493, -28879, -25035, -22961, -19754, -16625, -12869, -9065, 
    -4448, -100, 3168, 8255, 11160, 17599, 20521, 23802, 24648, 28467, 29127, 
    31098, 30623, 30104, 30488, 29579, 26659, 23564, 20621, 16923, 14035, 
    9867, 4671, 1350, -2973, -7181, -11314, -14697, -19138, -23323, -23906, 
    -28573, -29258, -31053, -30612, -29988, -29524, -28799, -26379, -24670, 
    -20703, -16224, -13369, -9042, -5023, -696, 3363, 7004, 11539, 16026, 
    20541, 22302, 24939, 25984, 29593, 31408, 30625, 29887, 30390, 28389, 
    26095, 23831, 20553, 17182, 14084, 7956, 4719, 1041, -3469, -8267, 
    -11213, -15751, -19183, -23418, -25063, -27260, -30433, -31141, -30366, 
    -31569, -30549, -28835, -26016, -24833, -21220, -18327, -15854, -10468, 
    -5053, -238, 3883, 7681, 10669, 14570, 18607, 22751, 25980, 26660, 29609, 
    31772, 30717, 32315, 31351, 28293, 27018, 24346, 20729, 17139, 15540, 
    9054, 4904, 476, -4253, -7437, -9793, -14133, -17612, -22426, -24263, 
    -28166, -27559, -29022, -30395, -32066, -30030, -28226, -28010, -24091, 
    -21949, -19437, -14262, -11264, -6919, -2115, 2161, 7634, 11195, 15161, 
    18305, 22454, 25184, 27140, 28902, 30743, 30805, 32215, 29441, 28924, 
    26448, 24040, 22025, 17829, 13453, 10917, 6231, 957, -3050, -7051, 
    -10086, -14760, -18592, -21299, -24494, -27049, -28842, -31939, -31019, 
    -31364, -29573, -30229, -26893, -23706, -22313, -19708, -13173, -10835, 
    -7911, -1860, 1254, 7202, 10619, 13366, 19346, 21818, 23558, 26309, 
    28906, 29601, 30980, 30908, 31406, 29834, 27388, 24300, 21147, 18855, 
    14201, 11197, 5781, 2450, -2804, -6815, -11535, -14548, -17408, -21868, 
    -23955, -26137, -27801, -28709, -30932, -31336, -30209, -28067, -27015, 
    -24878, -22151, -20103, -15586, -10847, -5265, -3233, 3118, 7487, 10381, 
    13887, 17180, 22599, 23592, 27685, 28954, 31079, 31828, 29331, 29975, 
    27761, 26054, 26489, 23364, 20026, 15397, 11267, 7949, 3785, -2107, 
    -5261, -9925, -15331, -17668, -22017, -23270, -27119, -29688, -31072, 
    -30062, -30300, -31107, -28303, -27397, -24663, -21886, -19986, -15057, 
    -10658, -7503, -3671, 1392, 5689, 10819, 14476, 19560, 21790, 22781, 
    27695, 27801, 29851, 32326, 30446, 31128, 28983, 27712, 25102, 21679, 
    20599, 16409, 11813, 8022, 2369, -1707, -5637, -9440, -13944, -17839, 
    -21083, -23468, -26592, -29778, -30000, -30938, -31568, -30705, -29990, 
    -28478, -25971, -21225, -19131, -15562, -12950, -7383, -3588, 908, 5510, 
    9556, 12697, 17980, 20561, 22201, 26817, 28565, 29728, 31126, 31395, 
    30382, 28134, 29036, 25698, 22174, 19942, 16744, 13761, 8266, 3119, 202, 
    -4778, -9966, -14181, -17752, -19892, -22503, -27499, -29088, -30241, 
    -30850, -31100, -30288, -29576, -27653, -26690, -22245, -20180, -16834, 
    -12353, -7826, -4467, 1742, 3741, 9098, 12205, 16883, 19110, 22943, 
    26619, 29574, 31237, 31252, 30769, 31316, 29293, 27164, 25417, 24162, 
    19697, 15876, 12883, 8307, 5554, 524, -5778, -10408, -12012, -15833, 
    -21301, -23929, -25840, -27255, -28988, -30020, -30916, -30258, -30181, 
    -28914, -26766, -23248, -19957, -15738, -13716, -9450, -5494, -1691, 
    3584, 8414, 12962, 17711, 18805, 23993, 26303, 28326, 30342, 30706, 
    29517, 30592, 29662, 28291, 26055, 23184, 19592, 16478, 13350, 8582, 
    3981, 795, -3950, -8625, -12390, -16577, -21491, -22729, -26977, -27562, 
    -30021, -30575, -31608, -30795, -29980, -27711, -26079, -22809, -20680, 
    -15933, -13936, -10244, -6543, -642, 4161, 7622, 10731, 18019, 19955, 
    23538, 26558, 26906, 30316, 30057, 31389, 31636, 29969, 28530, 27214, 
    23228, 20554, 17453, 13610, 9469, 4712, 726, -4354, -9600, -11568, 
    -15152, -19242, -22739, -25521, -28850, -29160, -30134, -29224, -31044, 
    -30508, -27408, -26647, -24322, -20288, -16598, -13403, -9628, -5769, 
    -1097, 3133, 8310, 13527, 15900, 19090, 21702, 25137, 27215, 27847, 
    29866, 31231, 30618, 28827, 27373, 26746, 23196, 19563, 18148, 15079, 
    9883, 5841, 928, -2907, -8855, -10998, -15555, -19872, -21494, -24565, 
    -27619, -29391, -29513, -30136, -30752, -29913, -28991, -27599, -25468, 
    -20756, -17232, -14375, -11051, -5497, -865, 2737, 7545, 10970, 15914, 
    17410, 20868, 25552, 27627, 29745, 29535, 30007, 29170, 30232, 28966, 
    26530, 22332, 21513, 18179, 14808, 11264, 5702, 3238, -2945, -7434, 
    -12258, -16200, -20217, -20861, -26266, -26460, -29238, -31200, -31406, 
    -30423, -28326, -29049, -26420, -23743, -21330, -19030, -13943, -9518, 
    -6920, -2142, 1712, 6923, 11181, 15061, 19062, 21628, 25859, 26969, 
    30316, 31513, 29881, 31045, 29174, 29314, 28069, 25161, 21430, 18718, 
    13212, 11308, 6964, 2786, -3109, -5993, -12495, -13476, -17426, -22574, 
    -24835, -27425, -29131, -30521, -30795, -30031, -29873, -27971, -26528, 
    -24377, -21971, -18971, -15042, -10714, -7224, -1225, 2313, 5615, 11070, 
    15495, 19160, 22128, 24448, 26039, 29040, 31418, 30787, 30553, 29816, 
    28264, 25622, 24540, 21187, 19427, 13540, 10866, 6619, 2874, -1296, 
    -7159, -11994, -13590, -18227, -22333, -25293, -27810, -28529, -30634, 
    -31420, -32105, -31532, -28877, -27852, -23516, -21466, -18010, -14572, 
    -9788, -6936, -2044, 1269, 6503, 10890, 13427, 18586, 20808, 23385, 
    26726, 28346, 29038, 30372, 31568, 30144, 29330, 26098, 25075, 22422, 
    18754, 15029, 12553, 8809, 2196, -2950, -4764, -10592, -13772, -17613, 
    -21882, -23838, -26161, -27440, -30788, -29418, -31692, -29979, -29305, 
    -27592, -24898, -21843, -18082, -15348, -11437, -8003, -2967, -304, 6306, 
    10777, 14735, 18820, 20621, 23516, 26734, 28953, 31084, 31241, 31091, 
    29451, 29333, 27619, 25211, 20889, 17677, 17224, 13057, 8019, 2916, -705, 
    -6602, -10375, -15083, -18788, -22120, -23681, -26812, -28384, -30624, 
    -29282, -32067, -30872, -28890, -27331, -25932, -23560, -19603, -15229, 
    -11626, -6576, -3524, 866, 4645, 8767, 15140, 16326, 19147, 22972, 25479, 
    28600, 30128, 30223, 31477, 31451, 30860, 28712, 26061, 23679, 19026, 
    16054, 12435, 6773, 2733, -1160, -5199, -9186, -12381, -16707, -20600, 
    -24161, -27418, -29180, -29121, -30561, -29846, -31406, -29789, -26986, 
    -25638, -23110, -21384, -16134, -12792, -7612, -3852, -278, 4835, 8041, 
    12899, 17800, 19587, 22929, 25644, 28081, 29703, 30475, 30784, 29405, 
    28977, 27290, 26118, 23163, 18595, 16897, 13233, 7563, 5882, 348, -5444, 
    -8186, -13911, -17066, -21174, -23944, -26411, -27822, -29870, -30566, 
    -29721, -30556, -29796, -29005, -25298, -22798, -21048, -16080, -12373, 
    -8892, -2663, -899, 4500, 8119, 13254, 16075, 19921, 23220, 26426, 27068, 
    28099, 29772, 30148, 31600, 28559, 28868, 25246, 22958, 19050, 18025, 
    11309, 10131, 4519, -225, -4088, -8265, -12818, -16908, -20794, -22776, 
    -25108, -27893, -31285, -29525, -30546, -30096, -31488, -27454, -25719, 
    -23491, -19814, -17247, -13170, -8840, -5444, -1730, 3175, 7269, 12978, 
    16079, 19055, 23238, 26068, 27221, 28890, 29689, 30936, 29961, 30032, 
    27082, 26194, 22561, 20047, 16862, 13426, 10220, 4289, 850, -2801, -8864, 
    -13540, -14882, -18183, -23711, -24485, -26935, -30884, -32324, -29382, 
    -32217, -30508, -28736, -26894, -23691, -19985, -17025, -12814, -9005, 
    -5903, -1525, 3591, 8265, 11598, 15579, 20536, 22391, 25803, 27048, 
    27649, 30708, 31419, 30353, 30166, 28418, 25929, 24844, 21468, 17723, 
    13498, 9472, 4737, 1903, -4202, -7303, -12072, -16139, -19104, -22225, 
    -24357, -26696, -30088, -29362, -31872, -29855, -31513, -28059, -26249, 
    -22992, -20991, -17055, -13187, -11179, -4852, -1726, 2776, 8155, 12464, 
    14629, 18295, 21987, 25561, 27928, 29260, 30707, 30742, 29974, 30190, 
    29827, 25916, 25560, 22281, 17675, 15032, 9325, 6412, 1648, -2558, -8290, 
    -11654, -14406, -18790, -23024, -25020, -28335, -29769, -30368, -30054, 
    -32487, -29624, -27222, -25105, -25999, -21744, -19148, -14737, -11135, 
    -6240, -1886, 4019, 6964, 11648, 14784, 18842, 22775, 25028, 27986, 
    29791, 28801, 30454, 31126, 29773, 28870, 26373, 23742, 20860, 19121, 
    14182, 10227, 5862, 2547, -2162, -6728, -11787, -15346, -17911, -22356, 
    -23520, -26129, -28219, -28730, -31204, -30219, -31267, -29554, -27888, 
    -23429, -23467, -19734, -15200, -10328, -5902, -1424, 3109, 6172, 11607, 
    13958, 18240, 21966, 24192, 27157, 28947, 30644, 31668, 31236, 30272, 
    29514, 27787, 23845, 20649, 18584, 13449, 10383, 5660, 2012, -1236, 
    -5969, -11303, -13774, -17628, -21900, -24027, -26970, -29351, -30453, 
    -30778, -32225, -30754, -27570, -26259, -24226, -23309, -20361, -14625, 
    -10603, -6062, -3799, 3228, 6742, 9135, 14393, 17513, 21461, 25370, 
    25932, 28454, 29919, 31740, 29831, 29696, 29932, 28094, 23795, 21731, 
    18317, 15423, 11778, 6459, 4518, -1554, -5485, -10000, -14107, -17093, 
    -21772, -25372, -25618, -29979, -29177, -30579, -29854, -30136, -28048, 
    -28422, -25977, -22052, -19232, -15046, -11319, -8937, -3672, 2148, 6639, 
    10005, 14599, 16138, 21972, 25025, 25540, 29943, 30160, 30169, 31187, 
    30811, 29265, 27108, 23938, 23586, 19949, 16068, 12115, 6344, 4044, 
    -1097, -6484, -8790, -14377, -17259, -19842, -22660, -27111, -27030, 
    -30287, -30151, -30206, -30379, -28976, -28699, -26590, -22560, -20734, 
    -16773, -10855, -8890, -3719, 328, 5648, 10085, 12461, 16756, 20545, 
    22587, 25723, 28469, 31091, 30132, 30903, 29300, 30000, 26614, 25772, 
    23453, 19570, 16938, 11821, 9414, 3001, -769, -6383, -10375, -14047, 
    -17407, -21247, -24945, -26874, -29137, -28830, -30373, -31888, -30809, 
    -28125, -28094, -24864, -22907, -20166, -17098, -12481, -8386, -4726, 
    -1197, 3859, 9039, 13706, 17704, 19258, 22952, 25910, 26914, 30055, 
    29819, 31176, 30606, 28216, 28005, 24371, 22001, 19846, 15540, 12782, 
    8604, 3422, 49, -5405, -8705, -12604, -16037, -21196, -24776, -26326, 
    -27891, -28772, -31663, -30398, -29028, -30124, -28144, -27307, -23600, 
    -20073, -15313, -13235, -9170, -5854, 469, 3577, 9907, 12649, 16738, 
    19835, 22966, 25891, 28546, 28757, 30767, 30300, 31307, 30530, 27502, 
    25597, 22678, 20242, 16585, 12704, 8838, 5469, 1629, -3953, -8111, 
    -12515, -16134, -19344, -22658, -25632, -27888, -29676, -30759, -29838, 
    -31044, -28771, -29141, -26330, -23599, -19840, -16297, -12722, -9766, 
    -5441, 1175, 4904, 8484, 13311, 16223, 19713, 22664, 26023, 27116, 29818, 
    30152, 31126, 31088, 29775, 28375, 25882, 24734, 20386, 17479, 12610, 
    8897, 5443, 1558, -4357, -7906, -12959, -17327, -19108, -22854, -24720, 
    -26739, -29410, -31560, -29833, -30790, -30648, -28846, -27499, -24628, 
    -21322, -17049, -12645, -9283, -4183, -236, 4704, 7499, 11116, 16134, 
    19283, 22435, 24993, 27603, 28972, 30116, 31537, 30633, 30691, 27417, 
    26520, 25495, 20993, 18618, 12171, 9978, 6912, 1593, -3385, -6943, 
    -11817, -16291, -19705, -21879, -24774, -26641, -29311, -31212, -32384, 
    -30941, -30639, -27512, -26748, -24283, -19421, -17090, -14943, -9771, 
    -6891, -2108, 2900, 6971, 11097, 14414, 18928, 21644, 24874, 27567, 
    30059, 29081, 31942, 30977, 30455, 30082, 26079, 24072, 20417, 17620, 
    14280, 10203, 6082, 456, -2746, -6689, -12030, -15426, -20306, -22774, 
    -26365, -27031, -28141, -30001, -31707, -31171, -28710, -29509, -26933, 
    -25207, -22297, -19583, -14519, -11285, -5293, -610, 2408, 7678, 12537, 
    14549, 19472, 20648, 25980, 27197, 28472, 30090, 30609, 30415, 29799, 
    28208, 25966, 24602, 22384, 18635, 13583, 10268, 7802, 3641, -2564, 
    -7010, -10960, -14507, -18896, -20679, -24120, -25473, -30164, -30040, 
    -31775, -30515, -29745, -27944, -27687, -25276, -21518, -17412, -15823, 
    -11322, -6000, -2537, 2783, 6382, 10610, 15212, 18230, 22327, 25123, 
    27189, 27148, 29221, 30184, 30658, 30063, 29734, 27685, 23444, 21851, 
    17855, 15631, 10852, 6067, 1608, -3127, -6357, -9660, -14512, -19344, 
    -21955, -25247, -26812, -28415, -28655, -31296, -30203, -30212, -28634, 
    -27411, -23854, -22976, -18619, -14915, -12528, -6518, -3630, 3090, 6105, 
    9230, 14952, 18214, 21471, 25031, 26168, 28743, 30729, 30106, 30834, 
    31682, 27675, 25766, 25043, 23424, 17660, 14729, 11475, 6817, 3880, 
    -1294, -4347, -9045, -14125, -17607, -21038, -23829, -25600, -27353, 
    -29710, -30570, -31159, -30596, -27926, -27668, -24624, -21904, -19845, 
    -15058, -11430, -6706, -2325, 2341, 4546, 10061, 14458, 19326, 20898, 
    23868, 27299, 29271, 30600, 30213, 30721, 30258, 30819, 27382, 24286, 
    22367, 20887, 15991, 12770, 7485, 2681, -978, -6800, -10406, -12596, 
    -17562, -20519, -22243, -27911, -29045, -30189, -31030, -30029, -28892, 
    -29861, -26461, -25313, -23079, -19129, -15584, -11014, -9061, -4307, 
    1395, 5331, 8835, 14443, 16867, 19866, 23683, 25023, 28750, 28763, 31906, 
    31549, 31574, 29776, 26805, 27211, 23992, 18740, 16105, 12415, 7149, 
    4094, -811, -4026, -8676, -13054, -18190, -20617, -23923, -24993, -29582, 
    -30547, -31424, -31261, -30127, -28864, -27483, -25390, -22655, -19479, 
    -16811, -12366, -7833, -4210, 480, 5453, 8661, 13060, 17028, 21421, 
    22841, 26257, 27750, 29192, 31063, 30499, 31141, 30596, 27943, 26548, 
    23683, 21002, 16648, 12267, 8440, 4343, -1714, -4052, -9455, -14662, 
    -16761, -18871, -22707, -25772, -27610, -30027, -30273, -30510, -29153, 
    -27877, -26575, -26470, -23510, -19320, -15699, -12674, -7780, -4730, 
    127, 5559, 7598, 12519, 16929, 19866, 23501, 24474, 29297, 29748, 31835, 
    30239, 32134, 29562, 29492, 27322, 23382, 19665, 17488, 11381, 9221, 
    4436, 578, -4107, -9641, -13018, -16423, -20020, -21843, -25667, -27547, 
    -30234, -30779, -31561, -30853, -29783, -27792, -27395, -23875, -20919, 
    -15631, -13402, -8419, -3196, -346, 4190, 9045, 11648, 17217, 20740, 
    23074, 25785, 26679, 29077, 30819, 30508, 31740, 30293, 27062, 27224, 
    24251, 20101, 17457, 12169, 9364, 4909, -777, -3424, -7669, -10779, 
    -16772, -19159, -22367, -24497, -27730, -29460, -30673, -30708, -30031, 
    -29312, -28880, -27535, -23940, -21809, -17207, -13401, -10146, -5816, 
    -925, 3192, 6403, 11547, 16652, 19520, 22673, 25924, 27690, 31060, 29876, 
    30860, 32283, 31161, 28440, 27643, 24678, 21224, 18442, 14398, 9226, 
    5887, 231, -2928, -8422, -11271, -16560, -18435, -23636, -25427, -26509, 
    -29174, -31970, -30771, -30642, -30708, -28615, -26737, -25163, -22244, 
    -17336, -14208, -9181, -5502, -1437, 2963, 8040, 12994, 14024, 18701, 
    23430, 23685, 27870, 29322, 30994, 30980, 30501, 29764, 29502, 26673, 
    23643, 22354, 17323, 14538, 9622, 6679, 1327, -3455, -7233, -12567, 
    -14977, -18947, -22401, -24701, -28880, -29330, -29846, -30323, -30539, 
    -30877, -28778, -25714, -24257, -21481, -18506, -14104, -10486, -6811, 
    -618, 2976, 7375, 9483, 15389, 19139, 22320, 24170, 26000, 28222, 28702, 
    30525, 29629, 30761, 28487, 27233, 25519, 21856, 18794, 14341, 11278, 
    6827, 3294, -2514, -5490, -11799, -15309, -18975, -22085, -23209, -26348, 
    -29988, -29203, -30915, -31958, -30253, -28864, -26956, -23180, -22308, 
    -19103, -14378, -10082, -6689, -3450, 1884, 6871, 10852, 15562, 18640, 
    21098, 24034, 27454, 28339, 29230, 30407, 29655, 29918, 28148, 27155, 
    24977, 23025, 18573, 15325, 9939, 6674, 3377, -1269, -5325, -9931, 
    -15539, -18513, -21167, -23027, -25896, -27598, -30616, -31159, -31125, 
    -30531, -29048, -26391, -24086, -22483, -17852, -16331, -10882, -6765, 
    -1783, 988, 6584, 10083, 14106, 17905, 21160, 23461, 27647, 28984, 28343, 
    31658, 30665, 30708, 29629, 28274, 26365, 22031, 19126, 16673, 12343, 
    7428, 1809, -314, -4814, -11208, -14935, -18473, -21490, -24422, -26932, 
    -27318, -30389, -31028, -31659, -30952, -29734, -26900, -24762, -22177, 
    -18690, -16821, -11797, -6734, -2049, 1392, 5808, 9862, 13337, 18139, 
    19845, 24068, 26069, 28272, 29519, 29919, 31826, 29321, 27805, 27494, 
    25687, 22563, 19678, 14571, 12874, 6871, 3933, -1799, -5296, -9460, 
    -13365, -18413, -21500, -23333, -25976, -28588, -28853, -30806, -31247, 
    -28948, -29661, -27088, -26190, -22205, -18699, -15967, -12904, -7918, 
    -2982, 685, 6196, 9773, 13910, 16300, 19874, 24354, 26244, 28545, 30546, 
    28870, 31829, 30283, 29457, 26840, 25141, 22791, 19312, 14678, 12448, 
    8181, 4375, -365, -5603, -9910, -13060, -18661, -21635, -24921, -25671, 
    -28724, -29444, -30536, -32156, -31002, -30326, -27995, -25069, -22725, 
    -19785, -17558, -11333, -9542, -4888, -1154, 6607, 10504, 13805, 17299, 
    20794, 22447, 25479, 27703, 31008, 29876, 30788, 30505, 30150, 27446, 
    25775, 23205, 21552, 14952, 11671, 8837, 3764, -1762, -4523, -8672, 
    -13057, -17062, -20493, -24524, -24884, -26942, -28544, -29930, -30815, 
    -30961, -29226, -26710, -26253, -22446, -19504, -18284, -13239, -9391, 
    -3852, -225, 5244, 9797, 12648, 16590, 19660, 24209, 25506, 27538, 29556, 
    30825, 31649, 30049, 29479, 28922, 25507, 24281, 20947, 17146, 13224, 
    8454, 3573, 776, -3767, -7748, -13858, -17907, -21183, -24116, -26757, 
    -26980, -31076, -30737, -31233, -29618, -29122, -27950, -26520, -24127, 
    -21798, -16901, -13196, -8843, -3942, 682, 5212, 7623, 11674, 15324, 
    19012, 21677, 27100, 27973, 28492, 30357, 31396, 30745, 28373, 30136, 
    26362, 23622, 22223, 18376, 14041, 8395, 4389, 1119, -5582, -9123, 
    -12873, -16060, -18748, -23965, -25890, -28508, -29650, -29845, -31671, 
    -29548, -28389, -28931, -26024, -23095, -21003, -18028, -12930, -10589, 
    -4610, -1523, 4002, 6990, 11235, 15541, 20756, 23513, 26134, 28613, 
    30079, 31569, 31220, 30427, 29760, 29546, 25685, 22363, 20067, 17766, 
    14498, 10852, 5612, 942, -3082, -7397, -11992, -16558, -19148, -22555, 
    -27072, -28750, -28911, -30404, -29320, -30416, -31252, -28028, -26656, 
    -25382, -21328, -17024, -13377, -11045, -6094, -436, 1968, 8425, 11746, 
    14914, 19553, 20823, 24719, 27831, 28462, 29707, 30629, 30313, 29055, 
    28924, 26286, 25242, 21193, 18699, 13509, 9711, 4682, 830, -4101, -8168, 
    -10088, -15838, -19876, -22829, -23733, -26544, -29549, -30074, -31258, 
    -30594, -29364, -30052, -26978, -23603, -21846, -18361, -14940, -10709, 
    -7515, -1940, 2515, 5927, 10232, 16548, 19057, 22465, 24350, 27227, 
    28347, 30458, 30812, 30204, 29417, 28799, 26703, 24643, 21224, 16997, 
    14791, 10048, 5545, 2532, -1112, -6102, -11583, -14519, -18274, -21428, 
    -25414, -26882, -28340, -31153, -29008, -31223, -30532, -28680, -27370, 
    -23834, -21389, -19526, -14399, -9475, -5459, -1790, 2095, 7684, 9991, 
    14957, 18501, 21833, 24414, 27810, 28185, 28898, 31681, 31018, 31262, 
    29285, 26470, 24966, 21882, 19698, 15161, 10232, 7181, 2969, -1886, 
    -6225, -10201, -13219, -18359, -21718, -23582, -26495, -28397, -29820, 
    -31849, -31036, -31541, -30185, -27895, -24418, -21997, -18717, -15885, 
    -10202, -8610, -2542, 1099, 5793, 10357, 14603, 16307, 21475, 26011, 
    27657, 30089, 28753, 30359, 30939, 29051, 28434, 29012, 25693, 22445, 
    18655, 15675, 10755, 7203, 1352, -2322, -6855, -10166, -14644, -16799, 
    -22080, -23966, -27145, -30476, -31110, -30681, -31371, -30353, -29065, 
    -26641, -24383, -21198, -19128, -15124, -11100, -8147, -3746, 641, 5721, 
    9560, 12970, 17071, 20293, 23665, 26831, 27879, 30089, 30857, 30871, 
    30931, 29854, 28466, 25358, 24323, 20009, 14759, 12835, 6916, 1928, 
    -2536, -4369, -8980, -14537, -16547, -20178, -23051, -26069, -28636, 
    -29413, -30357, -31977, -29062, -30808, -28264, -24580, -22248, -18205, 
    -15280, -12227, -6952, -2372, 822, 4768, 9062, 14244, 18650, 19695, 
    23741, 26009, 29638, 30109, 29933, 31588, 31229, 28459, 27135, 25021, 
    23475, 18749, 16444, 12673, 8113, 4589, -97, -4308, -9876, -12535, 
    -15727, -21650, -23912, -26353, -27790, -28315, -30083, -31184, -31523, 
    -28492, -27768, -25418, -23485, -18722, -16079, -12725, -8467, -3420, 
    440, 5012, 9619, 13359, 16251, 19533, 25441, 24620, 27291, 31261, 29691, 
    30398, 31062, 30687, 27170, 25427, 21776, 19446, 16703, 12703, 9386, 
    4691, -1248, -3820, -9455, -13781, -16407, -20101, -23376, -26410, 
    -28673, -29831, -31447, -32373, -29778, -28463, -27791, -25099, -23731, 
    -20951, -15047, -12452, -8011, -5737, 105, 4396, 8806, 12573, 15731, 
    19402, 22706, 24304, 29849, 29393, 30236, 30957, 31248, 29574, 27633, 
    25626, 24318, 19563, 16532, 12916, 9719, 4080, 413, -5662, -7229, -11609, 
    -16405, -20350, -23011, -25489, -26934, -29960, -29500, -31523, -31803, 
    -29840, -29178, -26092, -22324, -21116, -17053, -14101, -7870, -5862, 
    -980, 4832, 7777, 12344, 15356, 19437, 23130, 24149, 28134, 30602, 29633, 
    29234, 30552, 29851, 28799, 26937, 22583, 21430, 17040, 13364, 9668, 
    6054, 115, -3545, -7830, -13465, -17088, -19409, -23092, -25789, -28229, 
    -28323, -29551, -30489, -29486, -29804, -27863, -26549, -25492, -20068, 
    -17086, -12172, -9583, -4229, -916, 2294, 7818, 11380, 16169, 18700, 
    21658, 27072, 27046, 28721, 31146, 30119, 31236, 29780, 28236, 26705, 
    23798, 20429, 17948, 14255, 10083, 5968, 288, -2963, -6256, -10949, 
    -16147, -19036, -22891, -25332, -26894, -28575, -29486, -29397, -31229, 
    -29338, -29749, -25836, -24037, -20775, -18532, -15510, -10578, -6086, 
    -1232, 3688, 8352, 12068, 14448, 18885, 20475, 24344, 28753, 28943, 
    30566, 30493, 30505, 29756, 29994, 27119, 23448, 19869, 19491, 13573, 
    10388, 4670, 1311, -3625, -8550, -12518, -14435, -17397, -21448, -24939, 
    -27853, -27643, -29772, -29242, -30890, -29751, -27170, -26621, -24002, 
    -22430, -18893, -13931, -11024, -5382, -1834, 2360, 6416, 9870, 14997, 
    19793, 21188, 26290, 27050, 30178, 30253, 30957, 30909, 28726, 28026, 
    28016, 23914, 20153, 19931, 13972, 10208, 5906, 1466, -3736, -6346, 
    -10643, -13584, -18720, -20781, -24024, -26260, -28759, -28392, -31084, 
    -29699, -29693, -28346, -27767, -23384, -20836, -19287, -15325, -11439, 
    -8004, -2262, 1754, 7299, 11357, 14832, 20119, 22336, 24455, 26525, 
    30224, 31311, 31547, 30830, 29854, 29970, 26932, 25471, 21024, 18445, 
    15564, 10558, 7407, 2226, -2856, -6311, -11589, -16055, -18137, -21794, 
    -24637, -26491, -27788, -29899, -29890, -29501, -30422, -28997, -25472, 
    -24334, -20981, -18923, -15213, -10810, -6934, -3436, 1643, 5549, 9037, 
    13588, 17792, 22278, 23262, 26225, 28516, 29180, 30826, 30011, 30158, 
    29873, 26490, 24505, 23340, 19433, 15987, 12573, 7038, 3363, -1324, 
    -5651, -11308, -14003, -18150, -22634, -24362, -26644, -29187, -29648, 
    -30265, -30368, -29889, -29153, -26538, -24454, -20929, -17813, -15363, 
    -10986, -8401, -4054, 1352, 6302, 10086, 13703, 19508, 21564, 24546, 
    28104, 28392, 28157, 30342, 30737, 29078, 29056, 27661, 24915, 22608, 
    18884, 13889, 11880, 8464, 3382, -2132, -5030, -10648, -13617, -16385, 
    -21391, -23265, -26838, -27459, -29647, -29595, -30646, -30935, -29071, 
    -27182, -26073, -21458, -19979, -15720, -11892, -8001, -3321, 568, 5330, 
    10195, 14310, 18709, 20952, 23253, 27521, 29145, 30181, 30807, 30734, 
    30745, 29259, 28380, 25667, 23376, 19382, 17744, 11909, 6888, 5302, 325, 
    -4487, -7768, -13310, -17200, -21261, -23595, -26349, -27975, -29612, 
    -30866, -29437, -30519, -29525, -29224, -24635, -22571, -19638, -16500, 
    -13008, -8111, -4143, -337, 5498, 9674, 12408, 15817, 20876, 22092, 
    26546, 29261, 28955, 29758, 31153, 30204, 29191, 29458, 27299, 22067, 
    21319, 15324, 13408, 7350, 4470, -75, -5675, -8485, -13471, -16531, 
    -20624, -24104, -27060, -27457, -30162, -30662, -31493, -30817, -28689, 
    -27620, -24773, -24411, -20946, -16899, -13434, -8582, -3205, -484, 5545, 
    7700, 13243, 16611, 20423, 22382, 27353, 27227, 28850, 30365, 30437, 
    32209, 28375, 28346, 26309, 24299, 21391, 18467, 11229, 7553, 5036, 
    -1199, -4853, -8000, -13110, -16394, -21112, -24598, -25725, -28004, 
    -28752, -31017, -31230, -29427, -29231, -27640, -25783, -24746, -19325, 
    -16254, -12407, -9582, -4891, -1067, 3943, 7736, 13044, 16518, 19731, 
    22182, 25138, 27671, 28338, 30335, 29389, 30631, 30506, 27947, 26506, 
    22867, 20330, 16037, 13973, 9362, 4842, -332, -3857, -8054, -12826, 
    -16562, -20598, -23180, -26164, -28260, -29653, -30331, -30277, -31446, 
    -30335, -29480, -27014, -24722, -20213, -17568, -14210, -9082, -4534, 
    -684, 2226, 8865, 12313, 15492, 19923, 23658, 25800, 27605, 30155, 29770, 
    29902, 30168, 30767, 27464, 24642, 23795, 20419, 15768, 12597, 10367, 
    5093, 1499, -4095, -7389, -12421, -16414, -20299, -21773, -24732, -26740, 
    -29211, -30348, -32155, -30929, -29950, -26989, -25968, -25392, -21382, 
    -18005, -14137, -10562, -7191, -825, 4002, 8288, 13122, 16897, 18703, 
    22461, 26219, 27418, 29591, 30749, 31277, 30631, 29878, 28308, 26640, 
    23345, 20601, 17632, 14622, 8586, 3996, 2533, -2928, -6279, -10939, 
    -15359, -18739, -22393, -25432, -27585, -30681, -30007, -29709, -31695, 
    -29431, -28219, -26607, -24720, -20997, -19238, -14071, -9815, -6056, 
    -2163, 1759, 7242, 10071, 14202, 19060, 21906, 25148, 25858, 27556, 
    28657, 29929, 32108, 30164, 29798, 28362, 23395, 20796, 17788, 13727, 
    10549, 5462, 2775, -2224, -7673, -11093, -13727, -19823, -21966, -26345, 
    -27380, -30444, -29496, -29924, -29782, -30920, -27913, -26763, -24792, 
    -22276, -18865, -13300, -11392, -6078, -3266, 2107, 6687, 9925, 14146, 
    18029, 21380, 23890, 26180, 27632, 30246, 30282, 29954, 31131, 30216, 
    28915, 24956, 21860, 17906, 15205, 9761, 7886, 2127, -1851, -5218, 
    -10562, -14149, -18045, -21249, -24062, -27688, -28005, -28954, -30651, 
    -31323, -29386, -29044, -27418, -23973, -23091, -17885, -15383, -12482, 
    -7229, -1734, 1921, 6422, 9947, 12764, 18326, 19815, 24555, 26264, 28735, 
    28440, 31837, 30649, 30402, 29299, 26001, 25084, 23110, 18416, 16242, 
    11303, 6042, 1929, -1408, -4800, -9323, -13707, -17263, -20626, -24407, 
    -26734, -28716, -31564, -30858, -32084, -30383, -27921, -28861, -25086, 
    -21604, -18894, -14080, -10624, -7732, -3592, 916, 5650, 8780, 13680, 
    18084, 22576, 23936, 25734, 28951, 31077, 31318, 32199, 29974, 30270, 
    26309, 26927, 21307, 21050, 14864, 11268, 8040, 4049, -533, -5761, -9694, 
    -14067, -16873, -20267, -24512, -25149, -29484, -29623, -31636, -30491, 
    -29462, -28936, -27335, -24644, -24325, -18992, -16736, -11886, -7730, 
    -4025, 156, 4986, 9082, 14817, 17623, 20640, 24408, 24812, 28895, 28918, 
    30157, 31256, 30359, 29711, 28223, 24002, 22755, 21104, 16445, 10683, 
    7110, 3687, 337, -3982, -9101, -12652, -16006, -20780, -22574, -24437, 
    -28293, -29977, -31896, -29510, -30921, -28693, -27712, -25902, -21620, 
    -20616, -17601, -12320, -7637, -3592, 2005, 4104, 7993, 14073, 15991, 
    21761, 22934, 26599, 28756, 29253, 31779, 29753, 31978, 30260, 29310, 
    26750, 21875, 20659, 16415, 13396, 9242, 4988, 649, -5179, -8857, -13745, 
    -18174, -18536, -22285, -25939, -28377, -29408, -30328, -31217, -32055, 
    -29781, -27510, -27109, -23961, -19578, -16331, -12954, -8916, -5447, 
    -120, 4743, 8520, 12538, 16756, 18976, 22937, 25223, 26782, 28756, 30620, 
    29394, 30272, 29524, 27490, 26424, 24005, 21848, 17462, 11819, 7880, 
    5087, -84, -3675, -7902, -10914, -16988, -18934, -24118, -26364, -27341, 
    -29375, -31786, -31870, -29274, -29764, -28586, -25815, -24796, -18822, 
    -17557, -13892, -9501, -5342, 545, 3482, 9044, 11431, 15816, 20794, 
    22341, 26587, 28961, 28639, 29817, 31485, 31680, 29867, 27545, 24551, 
    24937, 21583, 17101, 12993, 10596, 4877, -601, -4441, -8670, -10751, 
    -17341, -19086, -22953, -25504, -26182, -29869, -30801, -31066, -30546, 
    -30094, -27972, -27532, -24160, -19371, -17320, -12760, -9442, -5362, 
    -696, 3473, 7879, 12399, 15919, 18730, 22521, 25832, 27112, 27916, 29263, 
    30448, 30279, 30227, 29652, 24994, 24968, 21353, 18070, 13660, 8922, 
    5680, 1305, -2849, -7914, -12397, -16261, -18188, -21719, -24692, -27163, 
    -29575, -28636, -31654, -31386, -29972, -26644, -25745, -23617, -21459, 
    -17211, -13401, -11182, -6827, -627, 2388, 7369, 11539, 15455, 18465, 
    21208, 25169, 28958, 29797, 30654, 30187, 30568, 29105, 29116, 27464, 
    23024, 20981, 16869, 13676, 9887, 7380, 1712, -3807, -5484, -10841, 
    -15340, -18653, -22219, -25761, -26313, -28472, -29451, -30435, -32147, 
    -30381, -29098, -25150, -23647, -20329, -17615, -13633, -10622, -5593, 
    -301, 1215, 7763, 10390, 16176, 18067, 22406, 25912, 27469, 28154, 30405, 
    30780, 30904, 30957, 29166, 26394, 23897, 21614, 19013, 15375, 8762, 
    6068, 2425, -2466, -7783, -10479, -14230, -18034, -20304, -26585, -27822, 
    -28973, -29161, -30726, -30543, -30871, -29780, -26526, -25371, -21940, 
    -17260, -12956, -11976, -7281, -2170, 960, 6444, 10916, 14891, 18747, 
    22497, 23967, 26086, 30442, 31510, 32224, 29783, 30732, 30008, 26790, 
    25575, 22408, 18836, 14645, 9908, 6763, 2909, -2380, -6432, -11900, 
    -16267, -16940, -20992, -24900, -27794, -29770, -30069, -30121, -30195, 
    -30688, -29172, -27623, -25023, -22253, -19111, -14905, -10096, -6067, 
    -1886, 2707, 6377, 9993, 14118, 17660, 21130, 24215, 26536, 29593, 29644, 
    29872, 29661, 28995, 29006, 28531, 25503, 22529, 17653, 14866, 10207, 
    6459, 1464, -1087, -6009, -10849, -13218, -17767, -21012, -24542, -25719, 
    -27950, -30698, -30152, -30220, -30406, -28980, -28428, -26384, -21966, 
    -19222, -16283, -10181, -8650, -3868, 1374, 4659, 8955, 14737, 17680, 
    19958, 25296, 27798, 27896, 29881, 30804, 30614, 29100, 28171, 27646, 
    26379, 22707, 20079, 15066, 11164, 7829, 3680, -1469, -5632, -9310, 
    -15205, -16104, -21003, -24674, -26707, -29361, -29737, -30843, -30882, 
    -30138, -29739, -27213, -26488, -22316, -19430, -16314, -13015, -8200, 
    -2427, 383, 5825, 9063, 12071, 17295, 20898, 23334, 26557, 27354, 29886, 
    30808, 31249, 31913, 29503, 26844, 25897, 24322, 20126, 17052, 13040, 
    7136, 3195, -234, -4346, -9628, -13096, -15981, -20703, -23127, -26706, 
    -28381, -30442, -31634, -31919, -30205, -28931, -26771, -25149, -23288, 
    -19128, -14629, -12334, -7334, -4146, 539, 5534, 8413, 12837, 17463, 
    20000, 22928, 24925, 29279, 29836, 29780, 31093, 32001, 27895, 28057, 
    25445, 24145, 19877, 16496, 12363, 6958, 2793, -247, -5069, -9056, 
    -13292, -16410, -20443, -24081, -27373, -27017, -30008, -30798, -31386, 
    -30319, -29282, -27533, -25244, -22342, -19208, -15562, -12118, -8591, 
    -6055, 127, 4847, 8092, 12749, 18300, 20294, 24372, 26025, 27563, 28233, 
    29108, 30551, 30834, 28824, 28391, 26674, 22192, 20440, 16851, 14525, 
    8957, 5847, -7, -3439, -8449, -12743, -15936, -21200, -22936, -26159, 
    -27317, -30785, -31209, -30801, -29262, -30056, -27004, -27668, -23311, 
    -20640, -15442, -13285, -7294, -5415, 310, 4598, 8125, 12520, 17215, 
    20795, 23958, 25205, 28674, 30856, 30544, 30371, 32001, 30576, 29179, 
    27544, 23244, 22151, 17535, 12839, 10087, 5353, 859, -2458, -7803, 
    -11394, -15717, -19296, -22757, -26315, -28129, -28653, -29080, -31053, 
    -30900, -30512, -29422, -26742, -24436, -19665, -17569, -12506, -10191, 
    -4115, -1576, 3165, 6808, 11966, 16259, 20600, 23535, 26011, 26473, 
    28122, 30694, 30618, 30098, 29288, 27076, 27640, 24304, 20402, 17156, 
    13763, 8000, 5494, 1407, -2322, -8131, -11498, -17270, -21022, -22049, 
    -24056, -26229, -29117, -30415, -30758, -31222, -29948, -28655, -27529, 
    -24346, -20957, -18548, -15152, -9864, -5814, -1757, 3469, 7364, 11431, 
    17360, 18590, 22080, 24612, 28999, 28316, 30563, 31135, 30261, 31312, 
    27990, 25198, 24867, 22344, 18210, 14989, 9878, 5807, 674, -4358, -6029, 
    -11579, -14850, -18866, -22450, -25380, -25736, -28880, -29066, -30905, 
    -31128, -30168, -28545, -26679, -24671, -22120, -18413, -15626, -10161, 
    -7728, -3542, 3934, 6593, 10774, 15095, 18499, 22335, 24807, 26493, 
    30099, 29069, 31476, 32179, 30077, 29401, 27279, 25057, 22324, 19615, 
    16081, 11606, 6244, 2373, -3779, -6248, -10623, -15546, -18786, -21379, 
    -24479, -26613, -29006, -29979, -30305, -30297, -28736, -28740, -26803, 
    -25337, -20051, -19569, -15174, -11310, -6496, -2184, 2573, 6352, 9791, 
    14269, 17920, 23347, 23403, 26931, 27566, 29688, 30393, 31176, 31065, 
    29453, 26380, 25220, 21503, 18502, 13093, 11465, 7849, 1607, -2365, 
    -5575, -10781, -15155, -17395, -20690, -25416, -27256, -27193, -30168, 
    -29266, -31237, -30187, -28500, -28026, -26197, -21674, -18470, -14870, 
    -11043, -6495, -1336, 2549, 5152, 10134, 13953, 18233, 22246, 24263, 
    26956, 28417, 31052, 30632, 30400, 29668, 29680, 27136, 25013, 21743, 
    17325, 14069, 11652, 9073, 2190, -2188, -6369, -10871, -15344, -18551, 
    -22238, -25409, -25642, -28035, -31272, -29888, -30212, -28591, -29056, 
    -27778, -25260, -22120, -19136, -14934, -10122, -7250, -2757, 1642, 6716, 
    10876, 14362, 16535, 19427, 22703, 27012, 28888, 28717, 29671, 31210, 
    29355, 29503, 25845, 23984, 20945, 18846, 15183, 11562, 7424, 4340, 
    -1776, -5295, -10047, -14119, -17351, -21968, -23853, -26777, -28462, 
    -29280, -31000, -31995, -31393, -28668, -26923, -27106, -22271, -19970, 
    -16489, -10557, -6881, -2353, 751, 6711, 9450, 13526, 18477, 21300, 
    24415, 26556, 29016, 30066, 31324, 30802, 30208, 28016, 26474, 25532, 
    23449, 18664, 15280, 12237, 8416, 3527, -527, -3957, -8112, -12292, 
    -15732, -21978, -24082, -25377, -27050, -29997, -31378, -32053, -31294, 
    -27905, -28588, -24598, -23451, -18530, -16000, -12366, -7972, -4202, 
    174, 4223, 7907, 13208, 17559, 21160, 23051, 24632, 29911, 29854, 29666, 
    31042, 30582, 29142, 28936, 26766, 24684, 20608, 16312, 12555, 8759, 
    4412, 269, -4434, -8213, -12682, -15228, -19762, -23928, -25955, -27929, 
    -30017, -31472, -30317, -31062, -29562, -27757, -25767, -22615, -20691, 
    -17724, -12777, -8400, -5882, -665, 5012, 8995, 12644, 16714, 18470, 
    24000, 25763, 26677, 29945, 31339, 31252, 30217, 30795, 28581, 25397, 
    22539, 20537, 17455, 12697, 8211, 5119, -176, -3385, -10344, -13966, 
    -16045, -19310, -22326, -24523, -27725, -29299, -29827, -29901, -29979, 
    -31292, -28565, -26779, -23577, -19188, -17479, -13690, -8165, -5706, 
    -2059, 4807, 7848, 11562, 16358, 20142, 22949, 25953, 28036, 29441, 
    30727, 32167, 30916, 31027, 28760, 26127, 24362, 20743, 16536, 13268, 
    9302, 4367, -263, -2164, -7248, -12786, -14670, -19369, -22531, -25761, 
    -26286, -28628, -31615, -32394, -32154, -30396, -27105, -28121, -25388, 
    -21240, -17984, -14046, -10908, -4572, -1380, 5181, 6518, 12654, 15554, 
    19973, 22862, 25379, 26895, 29861, 29345, 31642, 30914, 29792, 29610, 
    25176, 24327, 20556, 16775, 13900, 8772, 4214, 1523, -3838, -8044, 
    -12183, -15586, -19678, -22183, -25704, -28189, -27626, -30469, -31727, 
    -30031, -29094, -27740, -27982, -22867, -22226, -17492, -14400, -10346, 
    -6378, -2602, 3668, 8582, 11961, 14644, 18384, 23224, 27021, 28716, 
    28159, 29474, 31536, 30428, 28307, 29971, 27354, 25006, 22001, 17518, 
    13339, 9927, 6479, 1719, -2908, -7887, -11067, -14309, -19929, -21395, 
    -25986, -27235, -29040, -29663, -31816, -31174, -28604, -28819, -27754, 
    -25115, -22630, -18346, -14142, -10234, -5319, -2987, 2823, 5499, 12062, 
    15441, 18383, 20503, 25071, 26934, 28713, 29255, 30490, 30868, 29854, 
    28769, 25753, 25416, 21385, 18070, 14859, 11164, 4815, 2025, -2720, 
    -6735, -11679, -15895, -19201, -21554, -25270, -26421, -27965, -28791, 
    -29740, -31094, -31515, -30256, -26372, -25916, -20172, -16560, -15085, 
    -9845, -6696, -1632, 3257, 5220, 11446, 15116, 19068, 21694, 23961, 
    26483, 27613, 28971, 29837, 31647, 30373, 29852, 27551, 24140, 23690, 
    19116, 15648, 9583, 7380, 1497, -2270, -5252, -11974, -15070, -17826, 
    -22718, -24757, -27290, -28789, -30386, -30471, -29339, -31008, -27981, 
    -26799, -25166, -21897, -19139, -15795, -11290, -7408, -2682, 2013, 5916, 
    10921, 13196, 18389, 22409, 23864, 26015, 29488, 29048, 29312, 30370, 
    29966, 28812, 26890, 25830, 21526, 19752, 15151, 11860, 6526, 1842, -990, 
    -5110, -10179, -13756, -17805, -19520, -24465, -27551, -27621, -29497, 
    -29072, -30494, -29731, -28327, -27438, -23570, -21741, -19072, -14182, 
    -11803, -8024, -3447, 165, 6130, 9800, 14186, 17330, 21415, 25132, 26836, 
    28890, 29528, 30031, 30324, 30294, 28491, 27792, 25864, 22166, 19880, 
    17083, 11619, 8291, 2510, -2075, -5864, -9792, -13840, -17864, -20898, 
    -23883, -26954, -28245, -31002, -30289, -30150, -30011, -29848, -27657, 
    -25607, -23289, -19457, -14485, -12043, -7851, -2495, 230, 6678, 9370, 
    14167, 17834, 21077, 24507, 27763, 28093, 29039, 31170, 29977, 29558, 
    28744, 27704, 25609, 23573, 20141, 15416, 12940, 6960, 3087, -743, -4273, 
    -9577, -14301, -18733, -21705, -23113, -25872, -27469, -30456, -29783, 
    -30500, -30375, -28964, -27952, -25479, -24154, -19189, -15273, -13212, 
    -8248, -4297, 1137, 4282, 8115, 14115, 18224, 21468, 24400, 25325, 29157, 
    29153, 30050, 31455, 30582, 29287, 27781, 25803, 22980, 19469, 16807, 
    12599, 9668, 5183, -190, -5769, -9532, -12712, -15288, -21481, -22544, 
    -26334, -28171, -30409, -28861, -31134, -30328, -29947, -28653, -26599, 
    -24164, -20555, -15451, -12744, -8680, -2988, 500, 4165, 8113, 13283, 
    15980, 19852, 22306, 25131, 27440, 30416, 29485, 31002, 30938, 30153, 
    27144, 25308, 23036, 19878, 15887, 14816, 10010, 4132, -836, -3361, 
    -7677, -13056, -16402, -20349, -23022, -25737, -27563, -28067, -30280, 
    -30085, -29798, -30168, -29115, -26573, -24303, -21739, -16869, -12120, 
    -9053, -5514, -1682, 2995, 7322, 11845, 15828, 19373, 23001, 25547, 
    27960, 29899, 31072, 30358, 32007, 29701, 28279, 25188, 23868, 19150, 
    16729, 12518, 9733, 3524, 2203, -3671, -7008, -12657, -14735, -19312, 
    -22623, -24678, -27312, -28696, -30625, -31135, -30997, -29115, -27411, 
    -25983, -22281, -21484, -17657, -13503, -8684, -4690, -1718, 4380, 8907, 
    11079, 15949, 19786, 23094, 26160, 28215, 29890, 29912, 30157, 30062, 
    29909, 28379, 26477, 22428, 20488, 18820, 12806, 8845, 5926, -271, -2939, 
    -7419, -12923, -15342, -19084, -23608, -23580, -26666, -30362, -30695, 
    -30271, -31067, -30156, -30208, -26013, -24099, -20354, -17765, -12998, 
    -9612, -7194, -1143, 4753, 8673, 11140, 15124, 19349, 22255, 26019, 
    25791, 30558, 30234, 32559, 30201, 29532, 29635, 25520, 23016, 20334, 
    18121, 13332, 8862, 5057, 1104, -4312, -5852, -11111, -16144, -19403, 
    -22401, -25687, -27725, -28598, -30812, -31760, -30735, -29147, -28156, 
    -26546, -23095, -22480, -17175, -13798, -10700, -5676, -566, 2047, 7288, 
    12239, 15466, 18188, 22340, 25304, 27427, 29909, 29442, 31713, 32563, 
    30370, 29562, 28257, 25931, 20958, 17332, 15141, 9714, 6642, 318, -2587, 
    -6683, -10109, -16122, -16903, -21409, -22981, -27584, -29316, -30486, 
    -29739, -29879, -28828, -28123, -26699, -24154, -20301, -18498, -14582, 
    -11929, -7707, -1780, 1986, 6467, 9476, 14975, 19207, 22109, 24549, 
    26495, 29089, 28880, 30982, 31688, 29450, 30347, 27102, 25374, 23116, 
    18207, 13621, 12012, 7962, 1811, -2468, -5355, -11182, -14265, -17040, 
    -21900, -23460, -26527, -29186, -30536, -31077, -31331, -28410, -27616, 
    -25838, -23714, -22544, -20336, -15875, -9463, -6919, -2597, 2481, 6634, 
    10546, 15139, 16887, 21189, 23365, 26654, 29419, 30501, 30490, 30918, 
    30151, 30140, 27866, 26270, 22125, 19193, 14273, 11051, 8003, 3061, -400, 
    -5569, -11116, -12902, -19342, -21259, -24456, -26968, -29518, -29862, 
    -32131, -29623, -29219, -28543, -28964, -25238, -22451, -20853, -15226, 
    -10638, -7101, -3796, 876, 6010, 10175, 12510, 18599, 21616, 24553, 
    26115, 27003, 31115, 29756, 29112, 31481, 29480, 27595, 25650, 22877, 
    18425, 16846, 13651, 9357, 1942, -1864, -5824, -9530, -13727, -16705, 
    -20444, -23364, -25126, -29265, -30456, -30898, -31329, -29138, -30095, 
    -27330, -26020, -22843, -19891, -16496, -12503, -7911, -4938, 701, 7015, 
    8788, 13112, 16884, 21107, 24076, 24775, 28238, 29757, 29830, 30198, 
    30445, 29401, 28866, 26574, 23270, 20113, 16531, 11741, 7981, 3610, -281, 
    -5919, -8948, -14338, -16599, -22203, -23037, -26486, -28238, -29324, 
    -30015, -31172, -31177, -29890, -28126, -25852, -22799, -21554, -16291, 
    -13894, -8564, -4519, 455, 4680, 7356, 13324, 17568, 21382, 21951, 25023, 
    27898, 28733, 29131, 30862, 29782, 31042, 28319, 26293, 24374, 21021, 
    16287, 11851, 9661, 3565, -1111, -4198, -9469, -13006, -18009, -20072, 
    -22114, -24842, -28833, -28355, -30456, -31382, -31109, -29481, -28282, 
    -24525, -24274, -19811, -18104, -12442, -10064, -4511, -606, 5667, 7594, 
    11374, 16893, 18542, 22936, 26213, 27550, 28343, 30429, 31065, 29665, 
    28902, 28036, 27266, 22603, 21714, 15390, 11602, 7132, 3282, 200, -5000, 
    -9817, -12002, -16108, -18948, -23325, -26507, -26617, -31104, -31602, 
    -30456, -30889, -30635, -29576, -25631, -23629, -19548, -15841, -11788, 
    -8209, -5683, -1067, 2121, 7790, 12522, 15079, 18197, 23120, 26465, 
    28224, 28915, 29877, 30479, 30558, 30860, 26981, 26303, 22791, 21772, 
    16908, 14612, 9194, 3973, 957, -3286, -6875, -11700, -17128, -21163, 
    -22848, -24487, -26648, -30312, -29815, -31815, -31165, -28208, -28965, 
    -27262, -25045, -21188, -18634, -13727, -8449, -5321, -308, 3312, 7855, 
    12364, 15776, 19022, 23241, 25878, 26484, 28444, 30814, 30256, 31721, 
    31018, 29468, 26543, 23576, 20357, 17219, 13812, 9065, 5678, 2542, -2780, 
    -7408, -10980, -16771, -20821, -23466, -25617, -27233, -28975, -29172, 
    -31589, -30107, -30734, -28832, -26795, -23315, -21349, -17865, -14739, 
    -10147, -5180, -1945, 2683, 8066, 10762, 15349, 19146, 22074, 25398, 
    27495, 27519, 31812, 30445, 29224, 30683, 27864, 25624, 23660, 22119, 
    18352, 15078, 10604, 5894, 1903, -3504, -7204, -12004, -16057, -18054, 
    -21022, -25701, -27519, -28843, -29377, -30195, -30499, -28990, -28290, 
    -26148, -26008, -21752, -16838, -14650, -10750, -4360, -2228, 2697, 7326, 
    11678, 14964, 18187, 22960, 23255, 26512, 29898, 29786, 30781, 29005, 
    31640, 29503, 26693, 23716, 21235, 18457, 13744, 9278, 7422, 1933, -3403, 
    -5706, -11900, -16256, -18226, -22429, -24017, -27774, -29136, -29676, 
    -30815, -31769, -31161, -28564, -27838, -23613, -21126, -20138, -14131, 
    -10452, -8222, -2221, 2287, 6750, 10854, 14721, 18762, 22326, 24508, 
    26822, 28974, 30402, 31022, 30327, 30877, 30661, 25610, 23912, 21892, 
    19309, 15335, 11587, 6301, 1964, -453, -5563, -10439, -14332, -17999, 
    -21428, -24696, -26277, -29618, -29405, -30564, -32224, -30446, -27213, 
    -27594, -24347, -21211, -19590, -14626, -11510, -6681, -3002, 1305, 6949, 
    10224, 15064, 17842, 21065, 24845, 26086, 28742, 28834, 30764, 30086, 
    30390, 28877, 26811, 24828, 21359, 17745, 14986, 11182, 8392, 3303, 
    -1089, -6850, -10458, -14394, -19110, -21469, -24988, -26399, -28346, 
    -28992, -31595, -29811, -29525, -28380, -26928, -25281, -21581, -19561, 
    -14866, -12215, -7426, -3260, 594, 4841, 10460, 13814, 17005, 19875, 
    24989, 25524, 27358, 30856, 30741, 30548, 30930, 29009, 27589, 25963, 
    21728, 19957, 17198, 11193, 8571, 4571, -1911, -5658, -10973, -14384, 
    -17359, -20208, -23437, -26709, -27655, -29529, -31297, -29226, -30510, 
    -30189, -26743, -26708, -22717, -20013, -15663, -11074, -9357, -3246, 
    1569, 5495, 10810, 12450, 16713, 19945, 23254, 25017, 27413, 28744, 
    29740, 31041, 31110, 29318, 27166, 23750, 21721, 20310, 14291, 12988, 
    8295, 4326, -1025, -4819, -8574, -12688, -17360, -19753, -24677, -25127, 
    -28993, -30867, -30496, -30042, -31242, -28222, -29194, -25652, -23757, 
    -21393, -17396, -13405, -7604, -5300, -480, 4352, 8431, 14117, 15867, 
    21198, 23137, 27433, 28244, 29173, 30754, 30832, 29917, 30424, 27493, 
    26551, 23568, 20489, 16851, 12262, 7422, 5153, -151, -5708, -8990, 
    -13277, -16663, -19919, -23313, -27487, -28217, -28263, -30443, -30889, 
    -29821, -29141, -28384, -25367, -22654, -20317, -16046, -13170, -8766, 
    -5140, 1631, 5891, 8922, 11421, 16767, 20071, 22961, 24966, 29402, 30084, 
    31096, 31499, 30670, 30151, 27745, 24514, 23867, 20955, 15659, 12087, 
    7179, 5602, 544, -2439, -8087, -11900, -15648, -21652, -23280, -25469, 
    -26945, -28947, -30323, -30231, -31570, -29849, -28749, -25928, -24606, 
    -21273, -17226, -14154, -7758, -5043, -132, 2935, 7207, 12647, 17901, 
    18453, 22500, 25832, 27815, 28175, 31455, 31065, 30890, 29564, 28030, 
    26922, 23360, 19671, 17000, 14134, 8820, 5242, 1337, -3790, -8290, 
    -11934, -16230, -19326, -22713, -25558, -26886, -30294, -31061, -29569, 
    -31242, -28229, -28954, -26921, -23763, -21599, -17618, -14701, -9834, 
    -6101, -291, 2099, 6804, 13016, 15935, 18537, 23302, 24084, 26133, 27850, 
    30889, 31231, 31129, 28782, 28743, 27170, 22637, 20091, 17221, 13289, 
    9777, 5337, 1280, -3114, -8324, -13490, -17168, -18754, -22607, -26000, 
    -26608, -29604, -29906, -31293, -30658, -30483, -27642, -26798, -24276, 
    -20283, -18038, -14330, -10348, -4876, -2112, 2153, 7505, 12155, 15059, 
    19131, 22696, 25329, 28902, 30227, 31011, 32481, 29697, 30098, 27489, 
    27500, 25147, 21141, 17641, 15082, 9108, 5171, 1956, -3176, -7005, 
    -12723, -15694, -18762, -22379, -25371, -28509, -28505, -31034, -31203, 
    -31604, -29778, -29672, -26525, -22989, -21409, -17518, -14979, -11931, 
    -6072, -1518, 2926, 6186, 11612, 14404, 19260, 22850, 25291, 26615, 
    29458, 30004, 30632, 32447, 28948, 29103, 26322, 24125, 22283, 19503, 
    15734, 10468, 5636, 975, -2580, -7555, -11366, -15440, -18540, -21719, 
    -25757, -26836, -28143, -29453, -30948, -31126, -30128, -27592, -27957, 
    -25623, -20583, -17602, -14990, -11054, -6553, -2541, 2134, 6839, 9950, 
    14442, 19327, 21855, 24845, 27852, 29934, 29738, 30390, 31009, 29647, 
    28013, 26421, 24078, 20309, 18487, 14734, 11026, 8461, 2511, -2141, 
    -6825, -11176, -15451, -19618, -22964, -22854, -27288, -28748, -30346, 
    -31501, -30934, -29893, -28269, -26835, -24605, -22978, -17419, -15228, 
    -12282, -7040, -4145, 3344, 6808, 10966, 13180, 17920, 21832, 23148, 
    26809, 28011, 30742, 29277, 31020, 31501, 28943, 27160, 24795, 21192, 
    20073, 15290, 11242, 7176, 4006, -2011, -6399, -10831, -13252, -18630, 
    -20316, -23750, -26285, -27733, -30058, -29089, -29800, -29131, -29507, 
    -27628, -25953, -21017, -18945, -15958, -9976, -6824, -3049, 122, 5845, 
    10042, 13513, 17829, 20975, 23928, 26689, 28246, 28643, 30211, 31328, 
    29981, 30245, 27802, 26308, 22319, 19464, 14560, 12534, 6747, 3780, 
    -1241, -6685, -9125, -14241, -18045, -20667, -24363, -25722, -27991, 
    -30591, -31011, -30026, -29635, -30164, -27819, -26122, -21142, -19159, 
    -16171, -11307, -6718, -4837, 543, 6920, 11095, 14565, 17994, 20687, 
    23771, 27631, 28051, 29535, 30287, 31828, 29056, 28097, 28465, 25560, 
    23370, 17924, 16725, 12473, 7737, 4267, 234, -5385, -8667, -14392, 
    -17955, -20201, -24320, -26802, -29214, -29329, -31169, -30830, -29632, 
    -29108, -27884, -24315, -22483, -18216, -17274, -11138, -8617, -2507, 
    656, 4875, 8081, 14191, 16610, 20541, 23248, 25819, 29054, 29907, 30454, 
    31119, 29736, 27995, 26659, 26180, 23110, 19232, 16426, 13138, 9422, 
    3096, 1057, -4222, -10324, -12540, -16122, -20349, -22863, -26341, 
    -27430, -28674, -30744, -29951, -30646, -28549, -28204, -25571, -23221, 
    -20358, -15592, -14078, -7775, -4070, 237, 3754, 8753, 12933, 15693, 
    20548, 23955, 25699, 26616, 31038, 29148, 31436, 31735, 28553, 28915, 
    26445, 23488, 19781, 16690, 11459, 10469, 3138, -623, -4485, -10130, 
    -13470, -16279, -18969, -23029, -25172, -28671, -30627, -30233, -31605, 
    -31203, -28114, -28357, -24894, -23546, -19732, -16770, -14226, -8879, 
    -4321, 542, 4490, 7399, 13620, 17415, 20991, 23126, 24515, 28003, 29605, 
    29047, 31430, 30735, 30089, 28859, 26131, 23502, 21531, 17231, 12425, 
    9141, 4557, 1075, -3066, -8295, -12066, -15543, -21443, -22711, -25410, 
    -28115, -29913, -29744, -29634, -30785, -29165, -28884, -26854, -23273, 
    -21709, -15626, -14290, -9579, -5632, -340, 3749, 7642, 12695, 16002, 
    19829, 21363, 25492, 27319, 29176, 29750, 30137, 28799, 29100, 29525, 
    27086, 22317, 21158, 17805, 14573, 8827, 4159, 2211, -2600, -9037, 
    -10955, -15641, -19227, -23683, -26234, -28598, -28964, -29747, -31981, 
    -32295, -29851, -27677, -26811, -23836, -21902, -17357, -14104, -9763, 
    -6227, -978, 3995, 7818, 10488, 16433, 19328, 22092, 25293, 26598, 29844, 
    29656, 30459, 30685, 29770, 28252, 25524, 25791, 20088, 17186, 14441, 
    9512, 5912, 2102, -2627, -7234, -11436, -15179, -19407, -21692, -26019, 
    -28517, -28128, -30428, -31200, -31411, -30380, -28540, -25650, -22983, 
    -22614, -16436, -15151, -11599, -6423, -2236, 3577, 7241, 11303, 15661, 
    18613, 22789, 24284, 27246, 29017, 29330, 30487, 29934, 29705, 28290, 
    25240, 23325, 22389, 17495, 14421, 10382, 5720, 2308, -2930, -6714, 
    -10754, -16002, -20342, -22293, -24907, -27701, -29959, -31455, -29906, 
    -29758, -31006, -28832, -27527, -23572, -22561, -18765, -15884, -12300, 
    -7576, -3661, 1931, 6157, 11336, 14487, 19319, 21243, 24679, 26848, 
    29532, 30490, 31843, 29503, 28508, 30503, 26966, 24526, 20506, 18336, 
    14567, 10041, 6809, 3181, -1510, -5959, -9532, -14496, -18856, -22181, 
    -24018, -26003, -30409, -30345, -29757, -31064, -30483, -28994, -28366, 
    -25352, -20680, -17681, -13345, -10968, -5692, -2338, 2309, 5221, 9452, 
    13379, 19127, 21330, 24289, 27140, 29755, 30612, 30033, 30759, 30051, 
    30398, 27022, 23437, 21338, 20132, 13654, 10090, 7396, 1880, -2762, 
    -5680, -10014, -12804, -17956, -20183, -23188, -26250, -27972, -31001, 
    -30657, -30023, -30857, -28950, -28183, -25014, -22375, -19003, -14994, 
    -12037, -6904, -3839, 446, 6414, 9676, 13638, 18378, 20845, 25353, 25934, 
    26818, 30651, 31531, 29808, 30642, 28294, 27077, 24486, 21296, 19236, 
    15559, 12432, 7346, 3500, -899, -5220, -10869, -13047, -17511, -20939, 
    -23067, -27990, -27498, -29435, -30425, -30813, -29129, -28878, -28326, 
    -26435, -22916, -19969, -16039, -11724, -8437, -2616, -59, 5718, 9622, 
    14204, 16518, 22125, 23434, 26074, 29091, 28689, 31502, 30802, 30032, 
    29272, 27934, 25194, 21671, 20025, 17683, 12161, 8474, 4506, -753, -5270, 
    -8350, -13971, -19045, -19636, -23846, -27519, -28945, -29112, -30802, 
    -31105, -30780, -28536, -27284, -26150, -24365, -19699, -16129, -12150, 
    -9230, -3651, -56, 4724, 9787, 13785, 15819, 20836, 23041, 26398, 29282, 
    30581, 29920, 29620, 30275, 29037, 28622, 25603, 22157, 21251, 16367, 
    11379, 8558, 4830, -208, -5249, -7610, -11953, -15445, -20291, -24434, 
    -26205, -28267, -29570, -30330, -29881, -28811, -30943, -28616, -26515, 
    -21907, -20482, -17078, -12654, -9368, -3802, -158, 4268, 8782, 12520, 
    16828, 19529, 23618, 25813, 27603, 29003, 29689, 30102, 30225, 28447, 
    28907, 25566, 23603, 19402, 17663, 13060, 8451, 3945, -340, -5044, -7353, 
    -12230, -16164, -19505, -24096, -25656, -28525, -29161, -31319, -31853, 
    -29889, -31000, -27997, -26035, -23686, -19785, -17225, -13238, -8067, 
    -4729, -415, 3432, 7773, 13149, 15298, 19342, 22535, 24971, 27217, 28686, 
    30411, 30632, 31189, 30077, 27421, 25414, 22495, 21279, 16509, 14465, 
    9008, 4217, 1484, -5295, -8230, -13391, -14585, -17930, -22619, -25354, 
    -28141, -30167, -29807, -30992, -30478, -29886, -27975, -25728, -22549, 
    -22212, -17886, -14595, -9912, -4908, -2436, 3841, 6667, 11968, 14155, 
    18972, 23419, 25474, 27288, 28390, 31374, 29691, 30447, 30384, 29017, 
    28113, 24400, 21125, 18193, 13640, 11396, 6007, 480, -2345, -8172, 
    -11814, -16123, -18621, -20956, -24622, -27142, -28913, -29339, -31461, 
    -30365, -30480, -29871, -28198, -22698, -20842, -18683, -14786, -10205, 
    -5767, -2250, 3816, 7597, 10697, 15570, 20955, 22636, 26676, 27161, 
    27653, 30172, 30907, 31781, 28906, 28351, 25359, 25816, 20003, 18505, 
    15455, 9166, 6153, 2030, -3111, -7882, -12367, -16294, -18079, -22370, 
    -25130, -28052, -29644, -29950, -30169, -31113, -31329, -28109, -25529, 
    -24063, -21810, -17231, -14109, -9955, -6619, -1181, 3656, 6248, 10369, 
    14465, 19955, 22473, 25890, 26219, 29184, 30549, 30136, 32175, 29184, 
    29847, 27910, 24694, 21391, 18378, 13813, 10903, 5712, 1839, -1549, 
    -7131, -10507, -14230, -19193, -20459, -26050, -25622, -29756, -31259, 
    -30915, -31148, -30824, -28373, -26546, -24654, -20789, -18999, -14679, 
    -11907, -5923, -1620, 2682, 6020, 10531, 14867, 19722, 20534, 23920, 
    27101, 27148, 28393, 31207, 31384, 29479, 28366, 27388, 24652, 22382, 
    18638, 16150, 9954, 7484, 2516, -2274, -7342, -11743, -15048, -19357, 
    -20695, -23633, -26179, -28831, -30197, -29844, -31011, -31870, -27353, 
    -28198, -25345, -20766, -18554, -14645, -11244, -6924, -3338, 1626, 6447, 
    9952, 14691, 18479, 20012, 24284, 26801, 29966, 30274, 30086, 31262, 
    30510, 30153, 27585, 25079, 21896, 20067, 14964, 11938, 7215, 2492, 
    -1897, -4967, -8856, -13238, -18552, -19698, -22920, -26658, -28439, 
    -30887, -30573, -31344, -29532, -27991, -26269, -25430, -21162, -18167, 
    -14543, -12023, -8215, -4101, 627, 4734, 10692, 13329, 17123, 21996, 
    24193, 26697, 30140, 28731, 29650, 30751, 31032, 30573, 28615, 24378, 
    22587, 19112, 17160, 11277, 7643, 3865, -7, -6702, -8172, -13495, -18166, 
    -21929, -22705, -27169, -28535, -29770, -30609, -31359, -30277, -29911, 
    -28576, -24481, -22973, -19737, -16369, -13013, -6466, -4725, 663, 6517, 
    10049, 12951, 17248, 19235, 22512, 26550, 28012, 29567, 30644, 32019, 
    30702, 28280, 28093, 24652, 22529, 18642, 16561, 11900, 8737, 4205, -913, 
    -4397, -9699, -13143, -18376, -19926, -24351, -26536, -28243, -28380, 
    -29680, -29727, -30885, -30092, -27783, -26651, -22745, -21068, -17316, 
    -13449, -7388, -4858, 575, 5044, 9494, 11539, 16722, 20496, 23355, 27752, 
    29784, 28114, 29954, 30593, 30520, 29174, 27636, 26194, 21977, 18804, 
    16449, 12521, 7171, 3446, 1618, -4868, -9095, -12264, -15995, -21697, 
    -23554, -26117, -27106, -29154, -30725, -31796, -30882, -27880, -29147, 
    -26026, -22584, -20405, -15646, -11497, -8052, -5085, -543, 4576, 9529, 
    12909, 16440, 20034, 21722, 26337, 27541, 29713, 30019, 32172, 30849, 
    30442, 29192, 27327, 23810, 20981, 16641, 12770, 8894, 4443, 256, -3809, 
    -9891, -12647, -16433, -20255, -24009, -26322, -28784, -29766, -29763, 
    -32029, -31855, -28559, -28213, -27433, -23145, -21459, -17053, -12926, 
    -8840, -5654, 495, 2497, 7942, 12961, 16888, 19053, 23598, 26928, 27393, 
    28901, 30281, 32077, 30871, 29388, 28899, 25679, 23758, 21544, 17582, 
    13034, 10157, 5271, 72, -2979, -6985, -11404, -15031, -20040, -22385, 
    -25567, -27736, -29599, -29522, -31890, -29488, -29913, -27866, -26930, 
    -22964, -21432, -16235, -13050, -8387, -3710, -1223, 3937, 7285, 12606, 
    16136, 19459, 22846, 25056, 26596, 28922, 29835, 31100, 31465, 29809, 
    27991, 26783, 23487, 20687, 18110, 13810, 9111, 6593, 1225, -4533, -7608, 
    -12550, -15814, -21043, -22949, -25539, -27475, -28961, -32208, -31035, 
    -29391, -28718, -28663, -27773, -24074, -20898, -15911, -14155, -10668, 
    -6592, -292, 2932, 8279, 10815, 17100, 19077, 22281, 24012, 27103, 27709, 
    29541, 31466, 31757, 30437, 29587, 26879, 23746, 21034, 16627, 14555, 
    9175, 6874, 2573, -1961, -6080, -11865, -15745, -18975, -21580, -25300, 
    -26299, -28747, -28856, -30629, -30384, -29639, -29355, -27696, -24537, 
    -20574, -19073, -14229, -9260, -6731, -1921, 1911, 6603, 10767, 14852, 
    18048, 21247, 25931, 27260, 28648, 29811, 30332, 31015, 30332, 29160, 
    28318, 24801, 21891, 17597, 14011, 10233, 6833, 894, -658, -5738, -11389, 
    -14730, -19528, -21354, -25572, -26798, -28673, -29993, -29395, -31592, 
    -31326, -27912, -28077, -25034, -20507, -17862, -13709, -10945, -5625, 
    -2553, 1578, 6698, 9951, 14556, 18898, 22129, 26281, 26625, 29489, 29824, 
    30330, 32018, 31882, 29818, 27234, 24463, 22723, 18169, 15867, 11031, 
    5629, 1287, -2057, -6339, -9157, -14453, -18131, -21427, -23805, -26430, 
    -27921, -30691, -29838, -30302, -28503, -28853, -26080, -24304, -23643, 
    -17911, -16848, -11222, -7200, -2057, 1968, 5935, 11187, 13929, 18366, 
    20820, 23409, 26407, 28242, 30163, 30148, 32245, 29717, 29852, 27962, 
    25309, 22251, 17572, 16448, 11061, 8228, 1826, 87, -5566, -10769, -15740, 
    -17123, -21931, -25287, -26063, -30180, -30532, -29440, -31964, -30131, 
    -27746, -26723, -24775, -22401, -18463, -16096, -11117, -7785, -2790, 
    1044, 7435, 9827, 14372, 18152, 21998, 23725, 27470, 28597, 29116, 30207, 
    32105, 30200, 29253, 27801, 25905, 22911, 20260, 15233, 11986, 7013, 
    2985, -385, -6849, -10375, -14487, -16201, -21590, -23617, -25416, 
    -27756, -30757, -31742, -29594, -29439, -29230, -28242, -25075, -22637, 
    -20201, -15832, -11158, -7927, -3339, 622, 5213, 7664, 14120, 17721, 
    20858, 25012, 25921, 29319, 30165, 30058, 30993, 29654, 27973, 26568, 
    25131, 23150, 19076, 17120, 12726, 7610, 4920, 141, -4347, -9059, -13605, 
    -16971, -19714, -24449, -26737, -28972, -29917, -30739, -32242, -28878, 
    -28598, -29287, -24699, -23405, -19932, -15774, -13589, -9162, -4398, 
    2068, 3809, 8896, 12576, 16309, 21267, 22577, 27641, 26751, 29554, 31133, 
    30659, 30945, 27572, 27887, 26020, 22843, 18789, 16709, 11849, 7594, 
    4263, -174, -5343, -8439, -12125, -18237, -20613, -23056, -27327, -27708, 
    -29758, -28766, -29805, -30565, -28845, -28856, -27205, -24418, -19402, 
    -16235, -13452, -9326, -5394, 1515, 4391, 7799, 14138, 16409, 18497, 
    22684, 27340, 28487, 30568, 29292, 32232, 30450, 28502, 26400, 27456, 
    24353, 20252, 17084, 13348, 7726, 5982, -1017, -4539, -8667, -12298, 
    -15698, -19068, -23213, -26138, -27868, -27982, -29625, -30254, -31109, 
    -29055, -28638, -26426, -24260, -20946, -16117, -13443, -10007, -3587, 
    -1804, 3987, 7032, 12140, 15106, 20296, 22468, 26015, 27701, 28191, 
    30196, 30846, 29790, 28851, 27503, 27035, 23360, 19628, 17018, 12513, 
    9129, 5611, 1376, -3534, -8815, -11622, -15716, -19326, -21570, -25037, 
    -27516, -28974, -30256, -31243, -30519, -28821, -28090, -26171, -23002, 
    -21713, -17193, -12035, -8938, -5269, -1592, 3933, 8230, 11138, 16282, 
    18914, 22409, 24574, 27527, 28256, 29229, 29180, 29584, 30363, 27752, 
    25410, 24496, 20731, 19060, 14346, 9948, 4008, 1408, -3589, -7794, 
    -10907, -16529, -19598, -23605, -24718, -28750, -29763, -30364, -29153, 
    -29954, -31203, -29700, -25479, -25262, -21972, -17245, -13518, -10367, 
    -4440, -2383, 2309, 7955, 11811, 17102, 20931, 22751, 24774, 26051, 
    29161, 31729, 31117, 30511, 30386, 27825, 28164, 23442, 21626, 17712, 
    14562, 11270, 6104, 1938, -2748, -7658, -11154, -15223, -20360, -21203, 
    -24999, -28652, -27841, -30899, -30550, -31870, -30627, -29194, -27627, 
    -24354, -20303, -17269, -15138, -10655, -6668, -1009, 3355, 6763, 10921, 
    15374, 20257, 21399, 25766, 26127, 30345, 29993, 29042, 29964, 30804, 
    27473, 25869, 23514, 22105, 18204, 15097, 8929, 5544, 2452, -3181, -5771, 
    -10933, -15190, -17604, -21246, -25580, -28190, -29465, -31059, -31097, 
    -30976, -30421, -27605, -28294, -23827, -22858, -17506, -14203, -11546, 
    -6768, -1586, 3101, 8061, 12426, 14487, 17264, 21039, 24055, 27173, 
    28590, 30313, 29574, 31865, 29011, 29755, 28030, 24582, 20981, 19816, 
    15804, 10111, 7738, 2294, -3444, -6866, -10073, -14634, -19882, -22210, 
    -23438, -26077, -29298, -29674, -29930, -30904, -29753, -28284, -25548, 
    -24514, -22046, -19804, -13720, -10635, -7808, -1833, 1707, 6763, 8987, 
    14244, 18029, 22166, 24629, 28181, 27450, 29002, 30178, 30690, 29765, 
    29178, 26619, 25069, 20644, 18131, 15371, 10582, 7687, 3423, -962, -6460, 
    -11901, -13042, -19205, -22358, -24272, -26694, -29404, -29010, -30930, 
    -30299, -30456, -28569, -28408, -23727, -22324, -18796, -14893, -11722, 
    -7555, -3196, -223, 4676, 11558, 12895, 17505, 21464, 24386, 26321, 
    28707, 28751, 32250, 30021, 29357, 28566, 27110, 25443, 23389, 18485, 
    15653, 10327, 8170, 2949, -824, -5827, -10393, -14287, -16833, -20634, 
    -23365, -25226, -29573, -29358, -30840, -30747, -30779, -29412, -28944, 
    -24660, -23717, -18825, -15969, -12361, -8708, -3975, 1949, 5962, 8515, 
    12551, 17230, 21355, 24249, 26741, 27218, 29221, 30370, 29492, 30374, 
    30127, 26570, 27317, 23335, 19750, 15803, 13127, 8279, 4630, -1727, 
    -6106, -8948, -12687, -16526, -19974, -23850, -26256, -27865, -29925, 
    -31246, -31612, -31256, -29977, -27348, -26830, -23328, -20268, -17381, 
    -11301, -8270, -4591, 590, 4328, 7899, 12461, 17251, 19626, 23277, 26609, 
    28608, 28834, 30246, 30704, 28789, 29943, 26255, 26228, 23154, 20984, 
    15612, 12068, 8962, 4613, 81, -4816, -8510, -12619, -16326, -21419, 
    -24361, -25988, -27434, -30218, -31551, -31162, -31342, -28530, -28340, 
    -26738, -23158, -19936, -15716, -12549, -8756, -3621, -218, 2785, 9176, 
    13450, 15350, 19948, 22031, 25870, 27599, 29935, 29233, 30982, 31643, 
    29479, 28164, 27280, 23093, 21743, 16448, 13415, 8350, 3904, 558, -4523, 
    -7876, -11672, -16371, -18689, -24674, -25995, -26394, -29966, -30250, 
    -30146, -30444, -29633, -28324, -26781, -22852, -19765, -17616, -12425, 
    -8529, -4043, -20, 3778, 9519, 12184, 15517, 20551, 23487, 25883, 26674, 
    29887, 29395, 30255, 29554, 29084, 27205, 27225, 23104, 19968, 17807, 
    13373, 8295, 4798, 461, -4511, -6389, -13449, -15552, -20447, -22100, 
    -26110, -27569, -29527, -30557, -30010, -29414, -28546, -28326, -27148, 
    -24624, -22341, -17220, -14278, -10106, -6350, -334, 4615, 7637, 10457, 
    14521, 17917, 21836, 25588, 27047, 31114, 28723, 31604, 28969, 28798, 
    28168, 25234, 24515, 21055, 17260, 13228, 8710, 4878, 1885, -2645, -9118, 
    -11708, -14461, -20597, -23926, -25555, -27365, -28847, -29035, -31615, 
    -30600, -29121, -27957, -26005, -25019, -21127, -16866, -14602, -9507, 
    -6053, -1535, 2188, 7139, 10420, 15240, 17812, 21847, 24996, 28852, 
    29257, 31294, 29702, 31491, 30621, 29159, 27346, 23412, 21163, 17712, 
    14558, 9241, 6083, 2392, -1616, -7188, -11891, -14964, -17635, -21465, 
    -26524, -28448, -28838, -31916, -32475, -30600, -29135, -27649, -27908, 
    -24697, -20300, -17178, -14829, -9429, -5263, -2174, 2994, 5803, 11259, 
    16164, 18593, 20869, 24291, 26966, 30024, 29725, 31761, 30161, 30571, 
    27864, 27112, 24936, 21148, 18586, 13961, 10429, 5795, 2262, -4004, 
    -5309, -10415, -14399, -18956, -22894, -24616, -25708, -27416, -31100, 
    -30346, -31000, -29470, -29416, -27457, -23119, -22038, -19289, -14225, 
    -9563, -7268, -726, 3537, 5716, 11199, 14027, 17341, 21400, 24394, 27737, 
    28617, 29913, 31383, 30576, 29681, 29284, 26556, 25984, 22495, 18231, 
    14803, 10514, 6877, 3461, -1993, -6987, -11348, -13896, -16470, -22455, 
    -25046, -25730, -27684, -29220, -31146, -30159, -30127, -28420, -26467, 
    -23459, -22080, -17856, -14916, -11023, -5770, -1711, 1338, 5482, 10996, 
    13711, 17497, 21823, 25086, 28284, 27536, 30589, 30491, 30658, 28989, 
    29647, 27520, 24633, 20838, 17750, 15139, 11448, 7780, 4272, -2569, 
    -6073, -10551, -13561, -19092, -20656, -24354, -27887, -29111, -30207, 
    -32132, -31024, -30654, -28307, -28297, -26334, -21307, -19793, -15735, 
    -11526, -7648, -2855, 1565, 5490, 11095, 14366, 16521, 20235, 24606, 
    26406, 28641, 29573, 29697, 31068, 29850, 30954, 28316, 25208, 22327, 
    20473, 14590, 12793, 7737, 3110, -2662, -4046, -9441, -13970, -17676, 
    -21651, -23669, -25372, -26969, -30363, -30798, -31949, -29082, -29826, 
    -28804, -25952, -22265, -18827, -16273, -10784, -7611, -4130, 1807, 4984, 
    8298, 12516, 16434, 19759, 22649, 28074, 28612, 29573, 29824, 31511, 
    29873, 29742, 27707, 25354, 22546, 19273, 14914, 10937, 7546, 3847, 
    -1700, -6428, -7874, -12340, -16524, -21371, -23070, -26120, -29754, 
    -29323, -30405, -29656, -29155, -29682, -27179, -26205, -24225, -21035, 
    -15597, -12492, -8045, -3675, -312, 4417, 9449, 12458, 16347, 19743, 
    24792, 25278, 27529, 29875, 31028, 30446, 30060, 28707, 28378, 25949, 
    23852, 20338, 16184, 11443, 9913, 5053, -1052, -4118, -9169, -12773, 
    -16795, -19489, -22223, -25658, -26545, -29864, -30413, -30452, -30522, 
    -29561, -27587, -26132, -22636, -18423, -17263, -13204, -8254, -3902, 
    -30, 5433, 9644, 10914, 18133, 20091, 23164, 25856, 27243, 29207, 31395, 
    30151, 29765, 30344, 26326, 26932, 23058, 19798, 16383, 11744, 9542, 
    4342, -66, -3803, -8130, -11719, -15928, -20182, -23471, -25117, -28727, 
    -28479, -29089, -30844, -29152, -30088, -27657, -27255, -24579, -21274, 
    -15415, -13061, -9714, -4514, -172, 4487, 6890, 12294, 16066, 19276, 
    23218, 24553, 27329, 30077, 30919, 31559, 30911, 30099, 26967, 26531, 
    21956, 20683, 18286, 12532, 8055, 4153, 1596, -2497, -8706, -11147, 
    -17302, -17847, -21797, -24485, -28605, -29749, -30470, -31670, -29894, 
    -29192, -28872, -27782, -23927, -21030, -16298, -13406, -10185, -5687, 
    -1121, 3488, 8483, 12364, 15093, 19632, 23423, 24092, 28315, 29005, 
    31085, 30587, 30034, 28459, 29656, 25825, 23745, 20247, 16408, 13085, 
    10888, 5380, 1090, -3374, -7150, -10826, -17027, -18288, -22478, -24099, 
    -26544, -28171, -30442, -31346, -30365, -30644, -27973, -27051, -23603, 
    -19721, -17562, -12955, -9937, -5945, -990, 2483, 7778, 12544, 15627, 
    18566, 23581, 24697, 26656, 27647, 30092, 31443, 29315, 30924, 27298, 
    27003, 25099, 22070, 18470, 13899, 10140, 6361, 2688, -2949, -6758, 
    -10773, -16514, -19553, -22307, -24703, -27487, -29342, -30510, -31254, 
    -30585, -29772, -28315, -26521, -23379, -21045, -19101, -14141, -10709, 
    -6334, -2095, 1534, 7091, 10385, 15314, 18729, 21031, 24775, 26716, 
    29842, 29236, 30298, 31523, 29971, 28747, 27251, 25215, 20468, 17766, 
    14936, 9645, 5263, 2301, -2039, -7842, -12298, -16071, -18562, -22391, 
    -24084, -28251, -28868, -30684, -31902, -29514, -28812, -28358, -27400, 
    -25607, -21884, -18857, -14427, -11258, -7304, -2379, 2140, 7087, 10935, 
    14205, 18227, 21888, 24989, 26996, 28448, 31053, 29588, 30650, 31253, 
    28299, 27679, 24695, 23271, 19492, 13399, 10742, 5861, 2614, -1694, 
    -5947, -11715, -14830, -18174, -22000, -23922, -26681, -28680, -30606, 
    -31511, -29822, -29422, -28167, -26808, -25928, -21838, -18811, -15583, 
    -11172, -6082, -2879, 2340, 5402, 10427, 13639, 17887, 22663, 24097, 
    25314, 28610, 29185, 30425, 29207, 30710, 29066, 26252, 23903, 21668, 
    19916, 16560, 11118, 7297, 2479, -1532, -4170, -10121, -15047, -17295, 
    -20686, -23520, -25452, -28591, -29237, -30926, -29558, -29566, -28591, 
    -28015, -25825, -23518, -19807, -15944, -11277, -6198, -2044, 1023, 4483, 
    10555, 12643, 18283, 22482, 23994, 25431, 27802, 28867, 30371, 29815, 
    30083, 28981, 27683, 24752, 23678, 20067, 15232, 12902, 6943, 3304, 
    -2457, -6515, -10019, -13282, -16977, -20869, -23735, -26670, -28020, 
    -28915, -31211, -29848, -30608, -29011, -27860, -26227, -23595, -20749, 
    -14847, -12595, -6112, -4175, -160, 5367, 8969, 13624, 16291, 21229, 
    24584, 25722, 28413, 29984, 30432, 30168, 30539, 29607, 27613, 24221, 
    23016, 19485, 15065, 12795, 8616, 3299, -156, -3980, -8583, -11488, 
    -15374, -21202, -23625, -24968, -30194, -30171, -29841, -31419, -29345, 
    -29453, -27975, -25488, -23774, -20222, -17524, -11886, -9699, -5016, 
    720, 4822, 8687, 13929, 16714, 19115, 23951, 26773, 28465, 29121, 29923, 
    31136, 29718, 28926, 27373, 24869, 23811, 19226, 14873, 13065, 8938, 
    4836, -437, -3872, -8863, -13069, -16775, -20149, -23405, -26402, -27349, 
    -28984, -30918, -31607, -29943, -29291, -27049, -25636, -22833, -20553, 
    -17169, -13242, -8074, -3081, -963, 5633, 9561, 14416, 16185, 19690, 
    23930, 24902, 27402, 28825, 30536, 30762, 31890, 29199, 28848, 27389, 
    24062, 20472, 15588, 12630, 8446, 3842, -92, -3252, -8184, -13541, 
    -15850, -20032, -22070, -25035, -29219, -30067, -30660, -31570, -29183, 
    -28381, -29137, -25493, -22737, -20684, -16370, -12950, -8563, -5676, 
    -425, 3081, 7008, 12021, 15778, 20672, 23474, 24623, 27500, 30926, 30235, 
    29438, 30417, 30715, 28833, 26547, 23838, 20715, 17047, 13219, 8653, 
    5906, 682, -3676, -8376, -11174, -15442, -19910, -23263, -24741, -27848, 
    -29538, -30563, -32322, -29365, -28695, -29133, -27874, -23581, -19252, 
    -17918, -12030, -9706, -6204, -993, 3951, 7758, 13174, 15590, 19869, 
    21307, 25362, 27027, 29293, 30245, 30713, 30541, 30895, 28468, 26084, 
    23291, 21131, 18193, 13375, 10525, 4979, 2837, -5047, -7094, -12251, 
    -15673, -18661, -22211, -26480, -27023, -29186, -31605, -31261, -30343, 
    -28660, -27865, -25929, -24850, -22052, -18048, -13761, -9815, -4757, 
    -1029, 2336, 8191, 11779, 16663, 18635, 21929, 25176, 26498, 29359, 
    29916, 29947, 30885, 28750, 28580, 25909, 24072, 21790, 18735, 15567, 
    10568, 6273, 2844, -3842, -7078, -11547, -15205, -18549, -22284, -25810, 
    -27515, -29824, -28962, -30829, -29814, -29628, -30221, -26853, -25227, 
    -22763, -17666, -13858, -10177, -5854, -2732, 3502, 5215, 11396, 14607, 
    19056, 21740, 23987, 28644, 28262, 28851, 31642, 31645, 30777, 28412, 
    26310, 24428, 20279, 18355, 13392, 11936, 5953, 2128, -1538, -6495, 
    -10249, -14932, -17630, -20951, -24456, -26388, -29042, -28566, -30191, 
    -29923, -29253, -28158, -27530, -24816, -23039, -18500, -14503, -10972, 
    -4982, -1974, 647, 6674, 10004, 16083, 18659, 21861, 24388, 28153, 29523, 
    30515, 29346, 30692, 29177, 29717, 27783, 23521, 23440, 19365, 15219, 
    9830, 7229, 2404, -1852, -5292, -11000, -14380, -18154, -21484, -24902, 
    -26520, -29129, -29169, -30978, -30752, -30885, -28956, -27577, -25923, 
    -21982, -17811, -15523, -11556, -6768, -1955, 1715, 6276, 11509, 13971, 
    18276, 21046, 24185, 26215, 29974, 29796, 29792, 30781, 30111, 28692, 
    28441, 25277, 21684, 19097, 14875, 11360, 6834, 2477, -2664, -6215, 
    -9592, -14423, -18013, -19896, -23508, -27168, -28030, -30168, -31874, 
    -30112, -30128, -27548, -27305, -24598, -23607, -19114, -15764, -13177, 
    -6667, -2066, 1264, 6628, 11476, 12597, 17736, 19767, 24005, 27055, 
    29573, 31177, 29879, 30779, 28998, 30751, 28701, 24246, 23093, 19361, 
    16245, 12184, 8214, 2316, -2008, -4653, -8459, -12715, -18172, -21494, 
    -23550, -26700, -28234, -30192, -29497, -29676, -29111, -27961, -26215, 
    -25984, -21449, -20093, -16903, -12478, -8141, -2796, 484, 4862, 9595, 
    13588, 18871, 19926, 24703, 26244, 27095, 29499, 32061, 29986, 30016, 
    27887, 27715, 25966, 22877, 19818, 14650, 11513, 7035, 4720, -670, -4231, 
    -9344, -15157, -17030, -21005, -23485, -25783, -28710, -30067, -31469, 
    -31853, -31779, -30227, -27759, -25169, -24491, -20405, -16098, -10993, 
    -9212, -3360, -507, 4968, 10004, 12926, 18290, 20188, 24279, 25706, 
    27014, 29119, 32037, 31982, 30154, 28026, 27095, 26022, 22880, 20626, 
    16598, 13062, 9231, 2877, 565, -5679, -8343, -12855, -16880, -20124, 
    -23194, -25257, -26988, -30419, -31046, -31342, -31926, -29474, -29069, 
    -27400, -23313, -18332, -16577, -13507, -8957, -3661, 812, 4394, 7519, 
    13028, 17173, 20558, 22076, 26873, 28407, 29510, 31210, 30477, 29979, 
    29460, 28317, 27499, 23412, 20676, 18239, 11858, 9702, 4367, 1222, -3966, 
    -8968, -12056, -15343, -20257, -22931, -26412, -27608, -29798, -30867, 
    -32422, -30848, -29070, -28649, -26020, -22814, -21523, -15440, -13287, 
    -8641, -4856, -1249, 3484, 8353, 13005, 16991, 20632, 24452, 25296, 
    28907, 27902, 31179, 29694, 32244, 29811, 27687, 26831, 24281, 19261, 
    16376, 13640, 9399, 4163, -951, -3402, -6494, -12075, -16712, -19660, 
    -22765, -25938, -27705, -29067, -30240, -31744, -30223, -29027, -28741, 
    -27528, -24896, -19329, -17168, -12754, -9455, -6454, -592, 2732, 7599, 
    11999, 16640, 19311, 22750, 24201, 26254, 29202, 29687, 31180, 30309, 
    30580, 28323, 26407, 25363, 19177, 17041, 12959, 10533, 5701, 985, -2141, 
    -7839, -12887, -16562, -20771, -22498, -24949, -26395, -28562, -30409, 
    -30779, -31306, -30409, -28431, -26618, -25216, -21727, -18497, -13601, 
    -10739, -5898, -633, 3503, 7052, 12065, 14972, 19852, 21300, 24244, 
    27097, 28198, 29676, 31840, 31057, 29582, 28341, 27222, 22789, 21587, 
    18321, 13527, 9376, 4578, 2626, -2424, -7166, -11515, -16021, -20539, 
    -22084, -24919, -28849, -27628, -30596, -29284, -30723, -30518, -28932, 
    -26371, -24054, -20987, -17084, -15110, -8693, -6371, -1105, 2368, 7255, 
    10837, 14738, 18898, 22204, 26374, 28134, 28228, 30384, 31164, 30665, 
    30377, 29902, 26897, 26024, 22321, 19910, 13113, 9924, 6709, 2126, -3832, 
    -6715, -12528, -15113, -18727, -20570, -26007, -27497, -28572, -30354, 
    -30957, -30358, -30231, -29608, -25926, -24039, -21829, -18717, -12990, 
    -11122, -7622, -903, 2492, 6850, 9247, 14417, 18325, 21277, 24513, 27839, 
    28263, 29604, 30217, 30730, 29824, 28363, 26917, 23940, 23261, 18571, 
    15158, 9902, 5216, 1974, -2834, -7003, -9862, -16352, -18929, -21372, 
    -23956, -26498, -27459, -28509, -32049, -32170, -30160, -30338, -26099, 
    -24501, -21554, -19754, -14258, -9903, -6972, -3357, 1201, 7271, 9060, 
    15091, 17192, 22930, 24926, 28012, 28926, 29354, 30134, 30551, 30438, 
    28140, 27733, 24234, 21831, 18651, 14638, 11513, 7344, 2524, -613, -5292, 
    -9954, -15169, -18416, -20542, -24953, -25860, -28746, -30391, -31868, 
    -29620, -31182, -28525, -25795, -25997, -21759, -19184, -15640, -10307, 
    -6653, -4476, 369, 5288, 9905, 13226, 18732, 21561, 24326, 27032, 28325, 
    29375, 30126, 30626, 30861, 28945, 27247, 26307, 21418, 18813, 16488, 
    10347, 6470, 2792, -1656, -6207, -10640, -14185, -17893, -20770, -24050, 
    -27453, -29283, -30247, -30137, -30671, -31560, -30178, -28609, -25625, 
    -23022, -19536, -17477, -12220, -8027, -3096, 801, 4503, 9724, 14361, 
    17436, 21298, 24402, 26264, 29049, 29899, 28904, 29793, 31404, 29013, 
    28552, 24739, 23781, 19616, 16598, 11004, 8065, 2709, 782, -5617, -7770, 
    -14625, -16211, -20630, -22955, -25931, -30035, -31099, -30700, -30748, 
    -30412, -28486, -28541, -24480, -23989, -18526, -16723, -13220, -8219, 
    -5658, -11, 4977, 8604, 13262, 16738, 20280, 22535, 26240, 29125, 30020, 
    31423, 29699, 29391, 29796, 27732, 23936, 22939, 20943, 17323, 13079, 
    8507, 2969, -147, -4172, -8119, -12113, -15254, -19844, -23017, -25435, 
    -26878, -28144, -32078, -30877, -29675, -29470, -29225, -25873, -24810, 
    -20660, -15979, -12148, -8919, -6196, -882, 4032, 8256, 12454, 17063, 
    19725, 23424, 26256, 28066, 29458, 29898, 30975, 31500, 30446, 28404, 
    27034, 23825, 20850, 15284, 14149, 8390, 6314, 324, -5763, -7823, -12389, 
    -17574, -21152, -22613, -25647, -27178, -29573, -30204, -31058, -28822, 
    -29563, -28680, -26277, -23305, -20143, -15523, -13163, -10108, -5721, 
    -2087, 4357, 9045, 11132, 17012, 20852, 22995, 25413, 28503, 29864, 
    30955, 30886, 30642, 29606, 28538, 26257, 23545, 19773, 17850, 12284, 
    9820, 6673, 577, -4818, -8205, -12524, -16703, -19054, -22780, -25866, 
    -27968, -31222, -29382, -29943, -29763, -28658, -29800, -26165, -23271, 
    -21207, -17482, -14730, -8157, -4836, -1269, 2157, 6546, 13002, 15963, 
    21311, 22943, 27071, 27658, 29796, 29846, 32150, 30929, 30570, 28190, 
    25830, 23226, 20365, 16364, 13899, 9309, 6982, -655, -3230, -6840, 
    -11780, -15189, -20152, -21657, -23701, -27646, -30597, -30439, -30829, 
    -30568, -30033, -29945, -27769, -23830, -20065, -18833, -14652, -9969, 
    -6585, -1505, 4017, 7051, 12271, 14292, 18895, 23389, 25313, 27728, 
    28905, 30807, 29904, 29418, 30437, 28986, 27479, 23845, 21008, 17194, 
    13901, 9651, 5404, 1988, -2510, -6580, -11284, -15887, -17313, -23057, 
    -25942, -28466, -29704, -29074, -30652, -31352, -31028, -28525, -25513, 
    -24827, -22325, -18499, -13630, -10668, -6175, -2366, 2421, 7600, 10245, 
    15012, 18674, 22840, 25926, 28320, 29731, 29999, 29262, 30391, 30145, 
    29192, 27104, 23512, 20507, 17877, 14233, 11841, 6336, 2962, -2246, 
    -5652, -12264, -15689, -18755, -22159, -24904, -25883, -28668, -30225, 
    -28908, -30914, -29793, -29233, -26108, -24923, -22015, -17141, -15436, 
    -10653, -6440, -3113, 1351, 6617, 10051, 15236, 18240, 21543, 24115, 
    28091, 27328, 29082, 31309, 30016, 30418, 30010, 26509, 23983, 22296, 
    17775, 14715, 10427, 5678, 2771, -1006, -5705, -10856, -15294, -17345, 
    -20871, -23871, -25609, -27583, -29905, -31205, -29697, -30545, -29153, 
    -28311, -24085, -21921, -19407, -15909, -11756, -6599, -2512, 563, 6305, 
    8953, 14629, 17755, 20468, 24504, 27885, 29500, 28837, 30250, 31591, 
    31112, 29682, 27188, 25023, 22611, 20438, 15071, 11679, 8630, 1128, 
    -1604, -6768, -8978, -13897, -16781, -22281, -24142, -26160, -28889, 
    -28601, -30019, -31296, -29880, -27802, -28437, -24585, -23309, -19136, 
    -15740, -11946, -8978, -2995, 762, 6766, 9591, 13660, 17827, 19800, 
    25662, 27503, 27968, 30106, 31481, 31174, 30076, 30744, 27448, 24124, 
    21496, 19973, 14511, 12410, 8151, 3220, -1305, -4617, -10101, -14108, 
    -17408, -21721, -24219, -25230, -28524, -29627, -30579, -30840, -30806, 
    -28860, -28302, -24746, -23899, -18135, -16279, -12172, -8729, -3669, 
    534, 3525, 9368, 13312, 16928, 20851, 23588, 25919, 27358, 30330, 32204, 
    29931, 29302, 29286, 26885, 25443, 23608, 19939, 16670, 11342, 7632, 
    4114, -1958, -6120, -9724, -13725, -18102, -21622, -23385, -26523, 
    -28993, -30173, -30660, -31067, -30020, -28818, -28095, -26748, -22162, 
    -20124, -15816, -12038, -9306, -3524, 537, 5947, 8798, 14323, 16073, 
    21624, 22464, 24873, 27055, 31296, 30764, 32380, 30869, 29004, 26448, 
    26884, 22984, 18726, 16562, 12235, 10037, 3777, 775, -4273, -9610, 
    -13564, -16659, -19668, -23810, -25726, -29549, -30344, -29962, -29742, 
    -30957, -31350, -27527, -25506, -24054, -19389, -17994, -11791, -9272, 
    -3162, 1399, 4640, 7681, 12013, 15255, 19691, 21623, 26143, 27837, 28872, 
    29619, 32504, 30464, 31425, 28040, 26127, 24264, 19714, 16206, 12888, 
    8497, 6048, 487, -4228, -9227, -14087, -16544, -20730, -23426, -26089, 
    -28569, -29076, -30286, -30882, -30104, -29125, -27446, -27181, -24957, 
    -20973, -17417, -12856, -9012, -5109, -824, 4451, 8585, 13996, 15236, 
    20412, 23392, 24472, 28310, 29488, 30078, 32414, 31786, 29557, 29720, 
    26164, 22593, 21507, 18388, 13125, 9482, 5498, -456, -3179, -7348, 
    -12552, -16593, -20166, -22908, -25359, -26380, -30250, -30350, -29244, 
    -31026, -30835, -28064, -25404, -23206, -20567, -18756, -13016, -8248, 
    -4853, -249, 2546, 8181, 12672, 16868, 19388, 22966, 25244, 26687, 29204, 
    30437, 31362, 31322, 28242, 28218, 26755, 23862, 19350, 17984, 12562, 
    8806, 4853, 881, -3774, -8078, -12284, -16778, -20617, -23395, -24562, 
    -26642, -29869, -30817, -30296, -31643, -30385, -27675, -24664, -24391, 
    -19856, -17477, -13758, -9834, -5711, -2202, 2958, 5571, 11658, 16088, 
    19429, 23064, 24767, 27895, 29198, 31395, 31780, 31783, 29053, 28729, 
    27053, 25597, 19652, 18082, 15656, 9941, 4748, 1297, -2731, -5930, 
    -11048, -16678, -20147, -22791, -25636, -26560, -28974, -30093, -31798, 
    -29508, -29038, -27663, -27218, -24759, -20985, -18002, -14468, -10460, 
    -6986, -2031, 3398, 6259, 12882, 15891, 17871, 22826, 25044, 26907, 
    27469, 31270, 31209, 29781, 30245, 28948, 25808, 24558, 21004, 18379, 
    14899, 10717, 6607, 1729, -1347, -6421, -11315, -16357, -18379, -20279, 
    -25629, -27007, -29560, -30322, -31137, -29499, -30850, -30253, -26345, 
    -24254, -21487, -19281, -14926, -11250, -6178, -3231, 3013, 8126, 10928, 
    14498, 18679, 21776, 24736, 26538, 27544, 30455, 31246, 30256, 30112, 
    29849, 26894, 23871, 21896, 18679, 14343, 10945, 5306, 1485, -2852, 
    -6307, -9603, -15820, -19190, -21370, -23071, -27593, -29035, -30264, 
    -31204, -30637, -30812, -28959, -27273, -24503, -21390, -18373, -16315, 
    -11389, -7548, -3053, 1832, 4429, 10260, 14433, 16857, 21355, 25196, 
    27572, 29185, 29539, 30459, 31234, 29863, 28450, 28839, 24101, 22129, 
    19921, 15705, 11740, 8553, 1738, -2503, -5412, -9655, -12982, -18388, 
    -22023, -24818, -26092, -28774, -28372, -31207, -30850, -30686, -30613, 
    -27799, -25336, -23016, -18378, -16889, -9972, -5878, -1887, 1701, 5744, 
    10830, 13590, 17342, 22083, 24346, 26153, 28357, 28912, 30398, 31431, 
    30163, 29573, 27428, 25524, 23749, 20870, 15641, 10524, 7215, 2677, 
    -1485, -5342, -8867, -13804, -17095, -22426, -24235, -26162, -29533, 
    -30261, -31569, -30310, -30056, -29290, -26595, -23736, -23489, -19384, 
    -15913, -10320, -7659, -3434, 891, 5049, 8766, 15292, 16508, 22185, 
    25622, 26262, 28351, 29794, 31435, 31558, 29153, 29875, 27579, 26022, 
    21769, 20121, 16158, 11038, 9283, 4074, -1841, -4785, -8552, -11805, 
    -18180, -19860, -22616, -26069, -29330, -29426, -29617, -29415, -31491, 
    -29323, -26161, -24944, -23285, -19589, -16137, -13086, -8049, -3711, 
    -113, 4531, 8227, 12559, 16199, 21534, 23104, 26425, 29051, 28989, 30044, 
    31228, 31632, 30556, 29438, 24300, 21603, 19592, 17030, 11534, 9208, 
    3408, 33, -5034, -9110, -12769, -17284, -19574, -23890, -25434, -29541, 
    -29283, -31267, -31137, -30612, -29914, -28510, -26826, -21667, -20831, 
    -17034, -13748, -9145, -5765, 849, 4970, 7515, 12728, 17859, 19319, 
    23105, 25376, 27373, 30598, 29197, 31221, 30550, 28205, 27622, 24593, 
    23004, 19733, 15512, 11877, 9239, 5179, -17, -4314, -7654, -13284, 
    -15763, -20845, -23975, -24656, -27921, -28758, -30197, -30258, -29990, 
    -29671, -29362, -26128, -24258, -19023, -16312, -14218, -9581, -3841, 
    -1168, 2416, 8016, 12993, 16173, 20911, 24428, 25299, 28881, 30077, 
    30784, 29425, 30772, 30428, 29368, 27261, 22920, 22024, 17229, 14361, 
    9181, 6412, -577, -4266, -7775, -10876, -14649, -21044, -23943, -24847, 
    -27626, -29730, -30230, -30304, -30215, -29698, -28417, -25184, -23898, 
    -20367, -15775, -13503, -10163, -4898, -305, 3804, 9052, 12380, 15531, 
    18992, 21499, 24849, 27827, 28887, 31452, 29911, 31535, 30167, 27545, 
    26680, 23712, 21293, 17416, 14316, 9252, 6930, 652, -3319, -8405, -12682, 
    -14946, -18226, -22290, -26286, -27296, -29445, -31290, -31801, -31140, 
    -29387, -28412, -25543, -22786, -21094, -17989, -12515, -8321, -5955, 
    -1291, 3237, 8078, 11582, 16876, 18896, 22525, 25303, 27497, 29223, 
    29590, 30125, 29815, 30068, 27563, 26130, 23400, 20841, 18624, 13528, 
    10530, 5534, 1723, -2195, -6784, -11556, -14512, -20041, -23246, -25448, 
    -27185, -28929, -29456, -30744, -29748, -30466, -28861, -27873, -24038, 
    -20777, -17562, -15428, -10551, -6893, -562, 2454, 8170, 10370, 15705, 
    18772, 22495, 24571, 27061, 28253, 31850, 30927, 30950, 31391, 29107, 
    26956, 24834, 21835, 16801, 15713, 11020, 7392, 527, -2136, -5791, 
    -11262, -15148, -18159, -22234, -24137, -27985, -30240, -31088, -29215, 
    -30157, -29885, -29978, -26559, -25648, -22475, -18204, -14073, -12291, 
    -6237, -2817, 1685, 5587, 10326, 13202, 18387, 22314, 24308, 25411, 
    29383, 30018, 30596, 31618, 30188, 28769, 26923, 24971, 21927, 18038, 
    15657, 10956, 5626, 2270, -1668, -6210, -11341, -12693, -17581, -22931, 
    -23595, -26259, -30321, -30533, -30930, -30792, -30674, -29329, -26138, 
    -24669, -21732, -17227, -15554, -11337, -7165, -3097, 1668, 6001, 9348, 
    13285, 17769, 22214, 24889, 28398, 27747, 31831, 30001, 31423, 30508, 
    29957, 25896, 25024, 21151, 19790, 15084, 11776, 7151, 3158, -1625, 
    -5338, -11896, -12848, -17861, -21765, -22963, -27835, -28949, -29102, 
    -31447, -31470, -29951, -28678, -27124, -25759, -23275, -19675, -15924, 
    -12002, -6495, -4306, 1287, 5263, 11185, 13315, 17259, 20477, 23789, 
    26446, 28261, 31036, 29528, 30441, 29889, 29008, 29061, 24594, 23471, 
    18874, 14708, 10739, 7490, 2738, -948, -5747, -9125, -14467, -18122, 
    -20103, -22117, -26743, -29374, -29311, -30226, -31264, -30762, -29649, 
    -27895, -24949, -23183, -19912, -15184, -12311, -7483, -4148, 2520, 6612, 
    9249, 11831, 17122, 21420, 25132, 28022, 28210, 29460, 31329, 30136, 
    31584, 29955, 26359, 26965, 22271, 18929, 15538, 12534, 7844, 4098, -736, 
    -5146, -8875, -14702, -16760, -19435, -25006, -25391, -27803, -29555, 
    -29611, -30735, -31071, -29906, -27037, -24997, -24619, -20606, -15255, 
    -13005, -7848, -3923, -670, 6275, 10735, 11912, 16634, 21494, 23488, 
    26552, 28497, 29440, 29455, 31859, 29083, 29668, 27789, 26421, 22295, 
    19943, 17721, 13215, 8376, 3857, -1011, -4202, -9538, -12695, -17413, 
    -20948, -24005, -26139, -28632, -29030, -30344, -30757, -30722, -29502, 
    -28118, -25955, -22927, -21131, -16503, -13483, -9653, -6125, 1066, 3891, 
    9731, 12368, 16594, 20172, 22170, 25166, 28860, 29629, 30565, 30979, 
    30982, 29709, 26312, 26195, 24178, 20872, 16987, 14705, 8764, 4996, 77, 
    -3171, -8795, -13746, -16031, -19722, -21731, -25249, -29059, -29236, 
    -29573, -29900, -31129, -28002, -29421, -25948, -24266, -20026, -16700, 
    -12077, -10238, -4793, -980, 4646, 8432, 12095, 17467, 18693, 23835, 
    25950, 28437, 30069, 31419, 31883, 30922, 30217, 28291, 26739, 24040, 
    19838, 18086, 11660, 8285, 3944, 768, -2922, -8868, -10659, -17555, 
    -18883, -24145, -24847, -27522, -28176, -30965, -32001, -31554, -29884, 
    -27751, -26312, -23909, -19906, -16274, -12657, -9199, -5459, -1450, 
    5361, 6766, 11942, 17007, 18307, 22546, 26505, 27787, 28983, 30853, 
    31426, 31476, 29124, 29029, 25210, 24241, 19670, 18577, 12788, 9283, 
    4369, 1310, -2560, -8690, -12215, -16158, -20888, -22505, -25911, -26763, 
    -28680, -30060, -30902, -31698, -29044, -28567, -25583, -23901, -21193, 
    -18250, -14238, -10001, -4800, 233, 3467, 7090, 10310, 15216, 18054, 
    22549, 25733, 26522, 28800, 29621, 29085, 30626, 28686, 28650, 26100, 
    24234, 21301, 19365, 13107, 8515, 7177, 1401, -3350, -6240, -11867, 
    -14858, -19321, -22444, -25664, -25750, -29697, -29258, -30660, -30898, 
    -30679, -27429, -25597, -24005, -20213, -18943, -12715, -10435, -5729, 
    -2013, 3493, 6736, 11860, 14888, 19813, 21592, 25246, 28266, 30034, 
    29719, 30796, 29115, 29830, 28026, 26148, 24526, 22508, 17231, 14310, 
    11295, 7797, 2920, -3413, -5275, -11359, -16446, -18374, -23000, -25128, 
    -25674, -27793, -29962, -31266, -29762, -29015, -28887, -26445, -24762, 
    -21394, -18549, -14765, -9098, -7747, -1910, 3670, 5609, 10440, 15865, 
    17325, 20957, 24469, 27586, 28572, 29394, 30935, 31513, 31880, 30082, 
    25932, 26264, 21997, 18279, 13547, 10209, 6578, 2470, -707, -7004, -9837, 
    -14906, -17817, -21399, -25540, -26709, -28868, -31056, -32328, -30317, 
    -30165, -28907, -27735, -25256, -22724, -18672, -15298, -10421, -7452, 
    -1151, 1476, 7485, 10430, 14626, 17770, 21405, 23011, 27582, 29959, 
    29263, 30735, 31209, 29830, 28929, 27414, 24514, 22996, 19792, 15035, 
    11908, 7041, 2884, -2276, -6108, -8999, -12594, -17925, -22208, -23296, 
    -25259, -29248, -29785, -31422, -30853, -30803, -28881, -26436, -25205, 
    -21162, -18333, -16203, -12686, -7341, -2993, 624, 7211, 10668, 15041, 
    16215, 20586, 22571, 27801, 28219, 30213, 30956, 29944, 30587, 29627, 
    27079, 24364, 22771, 18801, 15926, 10946, 7823, 2846, -1004, -6716, 
    -10946, -12623, -17069, -19778, -24805, -25320, -28355, -28986, -30682, 
    -30927, -30361, -28758, -28851, -23675, -22382, -20232, -16438, -12086, 
    -7599, -4420, 95, 4627, 9255, 13400, 16215, 19670, 24468, 25290, 28885, 
    28871, 29883, 31547, 29832, 28580, 28044, 25464, 21078, 18245, 16947, 
    11722, 7726, 3524, 558, -5790, -8765, -13698, -17615, -20012, -22984, 
    -26960, -28287, -31167, -30313, -31064, -30097, -28417, -28047, -26056, 
    -23816, -19962, -16209, -11142, -8077, -2386, 161, 4398, 7880, 14033, 
    16892, 21719, 24726, 26823, 28789, 30052, 30586, 29404, 31172, 28423, 
    26399, 25486, 24250, 20971, 17014, 13007, 8353, 3065, -1121, -4245, 
    -8669, -13183, -16718, -19908, -22791, -26993, -28006, -29202, -30304, 
    -30964, -30717, -29547, -28454, -26242, -23459, -21016, -15792, -12079, 
    -8830, -4414, 156, 5644, 7895, 13340, 17018, 19864, 24238, 25645, 26467, 
    29597, 30173, 30319, 31767, 31069, 28183, 27021, 23525, 21304, 17069, 
    13360, 8461, 4197, 1537, -4913, -7948, -12622, -15127, -18637, -22593, 
    -25938, -29724, -30558, -28804, -30170, -30466, -30205, -28164, -26238, 
    -23291, -19150, -16801, -14557, -9195, -6675, -361, 4696, 7838, 10576, 
    16681, 19977, 22886, 24395, 26241, 29758, 31897, 31279, 30782, 30239, 
    28913, 24520, 23436, 19457, 17612, 14134, 9518, 5808, 11, -3240, -8362, 
    -14016, -16739, -19420, -23180, -25760, -28251, -29511, -30652, -31135, 
    -31505, -29619, -28943, -27097, -23521, -20286, -16149, -13893, -9288, 
    -3608, -917, 3166, 8244, 12281, 14545, 20088, 22907, 24483, 28217, 28812, 
    29560, 30708, 29585, 30735, 27642, 25759, 23041, 19909, 17673, 14189, 
    9088, 5688, 184, -3734, -8673, -10764, -15043, -18281, -21735, -26142, 
    -28033, -30402, -31143, -31144, -29258, -31514, -29231, -26168, -23096, 
    -21975, -18017, -13383, -8101, -3894, 72, 1983, 8199, 10990, 16332, 
    20421, 22028, 24714, 27501, 27717, 30302, 31450, 31459, 30303, 28852, 
    26157, 23915, 21515, 17207, 13865, 9294, 4735, 1931, -1915, -7346, 
    -12111, -15029, -20477, -23799, -25156, -27672, -28608, -29454, -30240, 
    -31404, -30408, -27349, -26494, -24614, -22557, -17118, -13768, -9883, 
    -6086, -818, 2655, 7239, 12027, 15569, 19363, 21697, 25248, 26553, 28466, 
    28323, 31615, 31101, 30139, 28317, 27318, 24014, 20748, 18987, 14570, 
    11175, 6794, 3435, -1713, -7702, -11750, -14762, -18574, -20713, -24269, 
    -26277, -28930, -30861, -29950, -30721, -29538, -29064, -25326, -24165, 
    -21073, -17456, -14873, -11528, -7751, -3076, 2255, 6758, 11231, 14680, 
    16660, 21197, 25255, 25658, 28105, 28643, 30491, 30878, 29393, 29579, 
    25934, 24683, 22217, 18352, 13996, 10529, 8281, 3082, -2294, -6068, 
    -11292, -14677, -19566, -21973, -24148, -28365, -29478, -30019, -30517, 
    -30884, -32034, -30399, -26429, -24984, -21572, -18526, -15758, -11870, 
    -7353, -1584, 1519, 7057, 11066, 14500, 18144, 21002, 23949, 26541, 
    27793, 29564, 32020, 31278, 28882, 28843, 27465, 25508, 23435, 19683, 
    16404, 10723, 8709, 2828, -886, -5658, -11225, -13719, -18090, -21999, 
    -24829, -27872, -29384, -29725, -30605, -31921, -30621, -30062, -27611, 
    -26319, -22349, -19487, -15386, -11724, -6597, -1944, 2720, 5829, 10983, 
    13006, 16591, 19822, 25043, 25739, 29714, 29912, 32232, 30640, 30437, 
    30474, 28231, 26455, 22430, 19360, 15200, 11727, 9059, 3278, -1940, 
    -5692, -10083, -11830, -18684, -21801, -24412, -27648, -29194, -29057, 
    -31327, -31730, -30895, -28763, -28197, -24444, -23144, -17996, -15693, 
    -10531, -7443, -3293, 1257, 5897, 8947, 13298, 18784, 20871, 23227, 
    26965, 29638, 29966, 29532, 30201, 29938, 28979, 28125, 25640, 22924, 
    19308, 15852, 12256, 7727, 4142, -1509, -4598, -8035, -14850, -17752, 
    -21972, -24109, -26365, -27888, -31429, -31095, -30011, -30327, -29016, 
    -29175, -25830, -23133, -19231, -15448, -11253, -7654, -2966, 58, 4954, 
    8315, 13590, 15689, 20157, 23180, 25743, 28388, 28010, 30610, 30900, 
    29282, 29359, 27288, 26327, 23469, 18698, 15557, 11418, 9599, 4174, 689, 
    -5650, -8981, -12696, -17072, -20070, -24014, -27322, -28143, -29823, 
    -30615, -30728, -30839, -29607, -28036, -25810, -23278, -20165, -16242, 
    -12170, -8494, -5511, 178, 4280, 8691, 12253, 16310, 21503, 23138, 26621, 
    27333, 30003, 30587, 31625, 30401, 28131, 28139, 25949, 23606, 20708, 
    17412, 11827, 9340, 4545, 368, -3645, -9559, -12448, -16451, -20139, 
    -23292, -26338, -28488, -29433, -30656, -31482, -30457, -28290, -27674, 
    -24661, -23336, -19556, -17323, -12763, -9313, -5029, -1305, 3336, 7935, 
    12413, 16917, 19979, 23225, 24904, 27216, 27670, 29616, 30871, 30718, 
    28817, 29113, 26032, 23691, 21290, 18819, 14463, 9235, 5867, 908, -3172, 
    -8042, -11672, -16553, -21328, -22758, -25400, -27602, -28018, -30248, 
    -30832, -31013, -28898, -28297, -26665, -25186, -20670, -18660, -14216, 
    -8432, -4870, -294, 3611, 7586, 12401, 16407, 19836, 21638, 24822, 28503, 
    28588, 29557, 31795, 29769, 29752, 29605, 26061, 22302, 20804, 16919, 
    14976, 9277, 4757, -192, -4322, -7916, -13046, -16398, -20610, -22143, 
    -25424, -27141, -29813, -31235, -30290, -30785, -29483, -27601, -26083, 
    -24976, -20880, -16756, -14638, -10367, -6760, -2340, 2263, 6135, 13257, 
    15673, 18908, 22017, 24184, 27307, 29404, 30162, 31241, 31487, 30845, 
    28600, 26599, 24819, 19575, 17404, 15063, 8480, 7390, 1894, -2500, -8326, 
    -10306, -15229, -19882, -23650, -25330, -27306, -28795, -29697, -30967, 
    -31211, -30361, -29181, -26625, -25195, -23134, -18405, -14426, -10198, 
    -6232, -2907, 2759, 7367, 10181, 16452, 17809, 20891, 25753, 28352, 
    29400, 28672, 29650, 30408, 30137, 28619, 28038, 24303, 22730, 19529, 
    13913, 11495, 5643, 2874, -2306, -6676, -11620, -14866, -19930, -20467, 
    -25486, -28699, -29389, -29230, -30695, -32458, -31022, -30084, -26428, 
    -23911, -22626, -18029, -14383, -11471, -6026, -1128, 1711, 4878, 10696, 
    15817, 16956, 21830, 22865, 26331, 29969, 30576, 30780, 30475, 29570, 
    29490, 26890, 24656, 21191, 18145, 14728, 11455, 7185, 3497, -822, -5592, 
    -10963, -12820, -18771, -22682, -23866, -26910, -28775, -29451, -29425, 
    -31384, -29431, -28252, -26863, -25865, -21193, -20204, -16248, -11548, 
    -6666, -4366, 2439, 4997, 11537, 15734, 17025, 19989, 25374, 27622, 
    29699, 30736, 29259, 30278, 30588, 29385, 27178, 24414, 22723, 18819, 
    15199, 11169, 6752, 3810, -536, -4834, -10526, -15352, -18271, -21503, 
    -24356, -25063, -28844, -30548, -31219, -29738, -29610, -30467, -28194, 
    -24909, -20790, -19882, -13983, -10763, -9177, -4056, 828, 4505, 10013, 
    12675, 16947, 21124, 22926, 26781, 28707, 29021, 30713, 31153, 29221, 
    29279, 27983, 25331, 22262, 19461, 14991, 10822, 7486, 4683, -1366, 
    -5350, -8588, -12114, -17612, -21965, -22224, -25495, -29182, -28577, 
    -31162, -31157, -30268, -29675, -27684, -25785, -21349, -18135, -16670, 
    -10400, -6622, -4571, 1811, 4809, 9071, 13986, 17283, 21266, 23546, 
    27272, 28591, 29883, 30578, 31184, 30129, 29137, 28029, 24927, 24209, 
    20593, 16913, 12658, 6801, 3027, -954, -4094, -9311, -13501, -17000, 
    -19785, -25065, -25777, -28353, -30694, -30001, -30892, -31399, -29463, 
    -27902, -25601, -23014, -20842, -17454, -11163, -9179, -3937, 366, 6177, 
    8256, 12942, 17240, 20882, 23695, 24792, 28014, 29819, 31310, 30384, 
    31013, 29441, 27812, 24082, 23436, 19603, 15948, 13535, 8969, 5959, 675, 
    -2946, -7693, -12664, -17938, -19509, -23675, -24975, -27567, -30062, 
    -29807, -31285, -31664, -30120, -28028, -26859, -23027, -20404, -15451, 
    -14061, -9440, -4198, -1031, 3448, 7799, 13825, 17071, 21066, 24525, 
    25060, 27513, 29572, 31887, 31497, 29860, 30300, 29327, 24458, 22738, 
    20048, 16923, 12521, 8060, 3677, 1799, -4500, -8102, -12165, -16241, 
    -20090, -23697, -26465, -27097, -29821, -30137, -30504, -30130, -30751, 
    -29226, -25728, -22817, -18745, -16774, -14040, -8452, -4802, 1218, 4573, 
    8324, 11866, 16087, 21191, 22338, 26180, 27999, 30331, 30437, 30593, 
    31693, 30072, 27501, 27342, 24524, 21044, 16749, 14128, 9296, 5969, 1142, 
    -2513, -8272, -12234, -14944, -20414, -23313, -25726, -27047, -30622, 
    -30512, -29286, -30449, -29934, -28880, -26051, -23928, -19706, -18524, 
    -13480, -9204, -4199, -818, 3958, 8139, 11511, 15995, 19949, 21909, 
    25747, 26830, 29445, 30272, 30517, 29578, 31256, 28376, 26204, 23968, 
    21706, 17237, 13583, 9055, 4393, -480, -3942, -7128, -11191, -16338, 
    -19457, -22512, -25812, -28609, -28366, -29479, -30360, -29968, -30750, 
    -28885, -24703, -24396, -19975, -18584, -14859, -10602, -5859, -923, 
    3933, 7795, 11211, 14075, 17854, 22111, 25548, 26982, 29221, 31817, 
    30511, 29850, 30382, 27941, 27895, 25001, 21233, 18022, 14623, 9431, 
    5876, 1009, -2869, -7260, -10210, -16434, -20827, -23145, -26094, -28042, 
    -29921, -30020, -30608, -30713, -30731, -28896, -26563, -23436, -21895, 
    -18069, -13854, -11639, -7258, -2083, 2666, 6408, 11032, 15259, 19278, 
    20484, 24099, 26328, 27782, 31836, 30909, 32133, 28762, 29308, 26753, 
    24710, 22386, 18684, 13783, 8937, 5584, 1984, -1567, -6225, -10832, 
    -15434, -18362, -21679, -23160, -28618, -30448, -29862, -31188, -31410, 
    -29812, -29774, -26957, -24627, -21476, -18463, -14341, -10231, -6844, 
    -1473, 1048, 7190, 10038, 14607, 18415, 21202, 24264, 27785, 28866, 
    29956, 31511, 30287, 31117, 30304, 26756, 24482, 20864, 18476, 15301, 
    10245, 7893, 1017, -2882, -5822, -10989, -13187, -19120, -21873, -25800, 
    -27796, -30090, -29795, -30653, -31666, -30987, -27802, -27619, -24065, 
    -22168, -19242, -14708, -10299, -7605, -3145, 1320, 5018, 9060, 14267, 
    17840, 23124, 24811, 27625, 27800, 30797, 29473, 30319, 30106, 29959, 
    28255, 25083, 21428, 19431, 16365, 11868, 7992, 2483, -1177, -6307, 
    -11256, -14799, -18293, -20738, -25778, -26241, -27830, -30792, -30232, 
    -30802, -31725, -28815, -27851, -24252, -23865, -17909, -14096, -11870, 
    -7524, -3966, 1301, 6556, 9060, 14674, 17387, 20967, 25116, 26583, 28099, 
    30081, 30312, 30915, 31173, 28728, 27807, 25162, 22414, 19272, 15201, 
    11044, 8002, 2180, -961, -4978, -9905, -13447, -17343, -20239, -23508, 
    -27655, -29415, -29691, -31790, -31043, -31418, -29792, -27872, -27096, 
    -22084, -20254, -17185, -13294, -8004, -3395, 1761, 5185, 9028, 15001, 
    18139, 19598, 25483, 24967, 28429, 29411, 31225, 30676, 30279, 28184, 
    27229, 25099, 23111, 19379, 16754, 13884, 9275, 3560, -1019, -4977, 
    -8180, -14467, -17376, -20055, -23120, -25425, -28596, -28954, -30486, 
    -29565, -31565, -28125, -28726, -25452, -23199, -19981, -16136, -13964, 
    -9169, -4011, -300, 5974, 9206, 13107, 18109, 20611, 23079, 26983, 28500, 
    31123, 29178, 30995, 31950, 28313, 28582, 24516, 22855, 20622, 16472, 
    12013, 10043, 4317, -417, -3176, -8274, -11349, -16866, -18596, -24121, 
    -24814, -27678, -29423, -31198, -30432, -30582, -29445, -28816, -26252, 
    -23233, -21599, -15786, -11697, -9558, -2807, 566, 3533, 8015, 12782, 
    17183, 20113, 22955, 25129, 28678, 28750, 30459, 30660, 29928, 28184, 
    28659, 27105, 23541, 20634, 16663, 13120, 10341, 3885, -1089, -5779, 
    -7918, -12751, -17662, -20339, -23261, -24751, -29446, -29399, -30486, 
    -29831, -28826, -28711, -26726, -27468, -22116, -19087, -16561, -12254, 
    -8223, -4367, 827, 4085, 8201, 13014, 15741, 19598, 23293, 24954, 29062, 
    30082, 30584, 31642, 32021, 30048, 28523, 27454, 23861, 22274, 17097, 
    12746, 8705, 4599, 742, -3578, -9034, -11689, -15924, -20318, -22728, 
    -25437, -27608, -28078, -30109, -30925, -30232, -30667, -28454, -26655, 
    -24820, -21687, -17318, -14062, -9280, -5346, -754, 4249, 8890, 12309, 
    14730, 20805, 21562, 26525, 28129, 29169, 30656, 30788, 31986, 31263, 
    28986, 24609, 22789, 20220, 16785, 12215, 9995, 6543, 1267, -4080, -7474, 
    -11583, -14919, -20213, -21316, -26665, -26877, -29495, -29656, -30065, 
    -30809, -28028, -27887, -26114, -25490, -21885, -18670, -14851, -9431, 
    -6677, -143, 4407, 6890, 12542, 15251, 18142, 22116, 24878, 26676, 30318, 
    31859, 30463, 31497, 29358, 29456, 25425, 24512, 22055, 19154, 14694, 
    9457, 5810, 2540, -1908, -6535, -10015, -14988, -17696, -23582, -24729, 
    -26631, -29450, -31359, -30667, -30953, -28723, -28593, -26845, -23169, 
    -22181, -17086, -14823, -11263, -6807, -3022, 4000, 7199, 10648, 13783, 
    19774, 21951, 23580, 27423, 28867, 29438, 31226, 30469, 30488, 28262, 
    26071, 25386, 22233, 19242, 14940, 11250, 5877, 2099, -2164, -5714, 
    -12146, -15651, -19609, -22281, -25328, -26410, -30120, -29770, -30400, 
    -30764, -29223, -27231, -26906, -26323, -21525, -18886, -14540, -11742, 
    -7091, -1383, 2231, 7789, 9261, 14397, 19642, 21212, 24475, 28275, 28388, 
    29567, 29828, 30572, 30195, 28316, 27999, 23735, 22190, 19577, 15793, 
    11525, 7108, 3490, -1531, -7430, -9619, -16263, -18672, -22097, -23947, 
    -26099, -29906, -31156, -30210, -31662, -31116, -28531, -26068, -24843, 
    -21684, -19786, -15193, -10652, -6003, -1154, 2149, 5253, 9387, 13296, 
    17577, 21579, 24720, 26787, 28248, 28753, 30351, 30414, 30612, 28687, 
    28201, 25261, 22774, 18339, 16939, 12102, 7439, 2996, -944, -6759, 
    -10495, -13271, -17347, -21104, -23628, -28508, -29322, -30566, -30235, 
    -30728, -28985, -29666, -27072, -24700, -22428, -17914, -15501, -9774, 
    -7447, -3656, 2583, 5833, 10352, 13939, 17557, 22204, 25009, 28001, 
    28178, 29716, 31524, 30014, 29974, 29287, 28372, 26610, 22010, 18426, 
    14865, 10341, 6461, 3049, -1282, -4936, -9403, -13488, -17189, -19923, 
    -24085, -24973, -29559, -30233, -32034, -31071, -31848, -28446, -27669, 
    -26732, -21088, -19586, -16850, -10645, -8166, -3099, 1249, 6778, 9280, 
    12550, 17706, 21016, 23691, 26545, 28474, 29547, 31054, 30865, 29122, 
    29258, 28090, 25650, 22099, 18548, 15944, 13792, 9024, 3824, -1441, 
    -3960, -8739, -12896, -18416, -19698, -22969, -26131, -27689, -29280, 
    -31603, -31310, -30649, -28098, -28673, -25361, -22317, -18319, -15329, 
    -12759, -7015, -3998, -664, 4433, 7840, 14231, 15334, 19395, 24008, 
    27126, 27760, 28790, 31407, 29700, 29773, 28739, 27170, 25426, 24269, 
    19363, 15972, 13560, 8906, 4032, -835, -5535, -9218, -12835, -17991, 
    -18622, -23437, -25163, -27883, -29481, -30331, -31087, -30366, -30873, 
    -26967, -25270, -23082, -19068, -15617, -12291, -8903, -4088, 1684, 3802, 
    8802, 13587, 17357, 18615, 23370, 25640, 28050, 28347, 29565, 29253, 
    30329, 30158, 27591, 25988, 23152, 21386, 16154, 13516, 8938, 5131, -398, 
    -4680, -8722, -11424, -16003, -20617, -22788, -25649, -27845, -29856, 
    -30934, -31224, -30129, -30186, -28413, -25551, -23385, -20156, -16216, 
    -12956, -9770, -4948, 964, 2340, 8223, 11826, 15219, 19676, 23507, 24816, 
    27652, 29801, 31549, 31050, 30942, 29323, 29055, 25430, 23973, 20428, 
    17243, 12405, 9541, 5327, -202, -3251, -9374, -11029, -16676, -19197, 
    -22949, -25223, -29072, -27531, -29959, -30500, -29120, -30477, -28235, 
    -25684, -23895, -20982, -16528, -12064, -9269, -5592, -1731, 2413, 6570, 
    11965, 15698, 20707, 22652, 26014, 27206, 29423, 31492, 31594, 30308, 
    31282, 27976, 26285, 22348, 20076, 17049, 12673, 10370, 6700, 2435, 
    -4528, -7643, -12588, -14324, -18803, -22017, -24962, -26199, -30815, 
    -30220, -30672, -29022, -30611, -28792, -26205, -24035, -20480, -16682, 
    -14327, -8375, -6291, -76, 1913, 5758, 11622, 14873, 17761, 20837, 24451, 
    27436, 29168, 31013, 29732, 31694, 28791, 29594, 25881, 24404, 20345, 
    19147, 15189, 9560, 6279, 2702, -2454, -8218, -10436, -16720, -19640, 
    -23786, -25680, -27944, -29958, -30408, -30321, -31161, -29141, -28686, 
    -25945, -22525, -21914, -17796, -13036, -9443, -5100, -1764, 1851, 7659, 
    10862, 14347, 18758, 20818, 25318, 26443, 29716, 30927, 29649, 29042, 
    28849, 28472, 27600, 23651, 21401, 17767, 13489, 10215, 6091, 886, -2438, 
    -7303, -10931, -14534, -18590, -20537, -24680, -28000, -28657, -30705, 
    -30867, -30235, -30062, -27922, -25611, -24225, -22581, -18874, -14555, 
    -10894, -6514, -1578, 1825, 6265, 11794, 15619, 18034, 20752, 24399, 
    26218, 28846, 30218, 31705, 31474, 30203, 29365, 26366, 24016, 20966, 
    19131, 14754, 10912, 5214, 2806, -1858, -5530, -10771, -15386, -18354, 
    -22966, -24676, -26947, -29396, -29207, -29419, -31851, -31570, -29639, 
    -27947, -24147, -21524, -20026, -14666, -12133, -7315, -1607, 2775, 4661, 
    9893, 13969, 17082, 21911, 23233, 27007, 29043, 28424, 30575, 30914, 
    29481, 28691, 28649, 25465, 20941, 17592, 15588, 11220, 6900, 2284, 
    -2118, -5829, -10750, -14249, -17669, -20633, -23752, -27428, -29018, 
    -30450, -29662, -29735, -28889, -28748, -26722, -24988, -21885, -18356, 
    -14281, -11153, -8147, -2778, 1451, 6227, 10119, 13222, 17564, 22326, 
    24316, 25077, 29066, 29484, 30381, 31459, 30751, 30542, 27278, 26627, 
    21913, 19894, 16182, 10947, 7715, 3933, -1785, -5929, -10584, -12940, 
    -17540, -20634, -25246, -25953, -28344, -29199, -29849, -30063, -29270, 
    -30197, -27310, -26011, -24012, -19931, -16214, -12371, -8105, -2726, 
    -19, 5368, 9489, 12828, 15819, 21607, 23896, 25555, 28644, 29536, 32137, 
    31578, 29320, 29122, 28231, 24996, 22974, 18383, 16504, 12750, 7577, 
    4640, 98, -4971, -8118, -12874, -16317, -20681, -24807, -26528, -26771, 
    -29677, -30774, -29655, -28578, -28847, -28877, -25994, -22973, -21110, 
    -16604, -13533, -9512, -3853, 1327, 4948, 8340, 13905, 16287, 19430, 
    23707, 27547, 28798, 29519, 30425, 31138, 30019, 29617, 28368, 24414, 
    23016, 18198, 17829, 12629, 7658, 3735, 197, -4774, -8704, -14133, 
    -16892, -19589, -23180, -25662, -27038, -30299, -30557, -31559, -31155, 
    -30663, -28437, -26685, -24013, -19533, -18191, -12578, -7635, -4381, 
    -1570, 4115, 7487, 13095, 15315, 19383, 22785, 26295, 27777, 29763, 
    30962, 30118, 30052, 29666, 29599, 24579, 23484, 19224, 16026, 13229, 
    7762, 4881, 182, -5734, -7895, -11139, -16917, -20491, -23956, -25022, 
    -26904, -28346, -29703, -30042, -31260, -29666, -27332, -27013, -23539, 
    -19740, -16893, -13026, -10057, -5452, -2161, 3095, 8776, 13477, 15565, 
    20657, 24343, 24545, 28189, 29959, 30757, 30765, 30468, 31482, 27290, 
    25615, 24798, 20920, 17651, 13358, 9094, 3891, 35, -5182, -9580, -12139, 
    -16984, -20908, -22072, -25177, -28784, -28990, -28817, -31035, -30020, 
    -30098, -28481, -27507, -23613, -19868, -17990, -14299, -9865, -5085, 
    123, 3643, 7397, 11623, 16610, 18981, 22740, 25933, 28087, 28625, 30815, 
    31465, 29687, 30128, 29291, 26329, 24249, 20805, 16710, 14497, 8740, 
    5192, 515, -3985, -7691, -12534, -15693, -20826, -21958, -25639, -28493, 
    -29552, -28785, -30317, -29507, -30192, -28300, -25486, -25565, -20185, 
    -15898, -14205, -9878, -6251, -2727, 3172, 7019, 11409, 14776, 18708, 
    22979, 25963, 27111, 27915, 28927, 29873, 30145, 28544, 29788, 27801, 
    25063, 22195, 17574, 15171, 9225, 4776, 1311, -3924, -7260, -9478, 
    -16859, -17624, -23129, -25393, -25872, -29508, -29477, -31054, -31212, 
    -29732, -28517, -28216, -24084, -22428, -19113, -13837, -10416, -5989, 
    -1231, 1979, 7228, 10136, 14143, 19188, 22809, 23861, 26330, 30173, 
    29463, 29403, 30812, 30699, 29274, 26795, 23604, 22012, 16577, 14538, 
    10075, 5707, 2579, -1656, -7096, -11180, -15833, -19018, -21808, -25865, 
    -26157, -29319, -28941, -30722, -31112, -30365, -29057, -27697, -25119, 
    -21806, -19268, -15185, -11174, -6367, -1146, 2242, 6039, 11330, 15689, 
    18094, 21553, 26170, 25634, 30113, 29363, 29729, 30947, 30361, 28822, 
    28077, 23288, 21415, 18149, 15511, 10569, 5928, 2086, -2614, -6269, 
    -9726, -13525, -19514, -22743, -24637, -28249, -27807, -30862, -29906, 
    -30764, -28580, -29178, -26459, -23455, -22857, -19023, -13419, -11629, 
    -6528, -2245, 2631, 7742, 9908, 13732, 18208, 22602, 24601, 26501, 29844, 
    30836, 30369, 29413, 30498, 29652, 27158, 24710, 22365, 17376, 13779, 
    12009, 8897, 3567, -2346, -5248, -10769, -15341, -18212, -20450, -25228, 
    -27063, -27783, -29182, -29905, -31400, -30588, -29096, -26909, -25472, 
    -22720, -19569, -14902, -11930, -6858, -2860, 190, 4999, 9841, 13238, 
    18120, 21840, 23924, 26466, 28123, 28325, 31864, 29393, 29137, 30306, 
    27462, 26925, 21747, 19044, 17436, 11710, 8489, 3182, -1381, -5587, 
    -9279, -13141, -17624, -21705, -24005, -26095, -28565, -30123, -30838, 
    -30452, -30737, -30154, -28968, -25749, -22117, -20332, -16832, -12354, 
    -7817, -2969, -459, 5166, 10283, 13629, 18032, 20840, 22736, 26741, 
    28575, 29955, 30621, 30915, 30006, 29151, 27908, 26315, 22501, 21181, 
    15596, 12077, 6437, 2712, 806, -4249, -8537, -12371, -17160, -19979, 
    -22871, -27122, -28698, -28070, -30244, -30221, -31239, -29645, -28148, 
    -26903, -23214, -19123, -16523, -13206, -7310, -3872, 196, 3634, 10612, 
    13484, 17267, 20124, 22876, 25720, 27989, 29926, 30781, 32649, 29374, 
    28339, 27477, 26622, 22875, 19517, 16490, 11685, 9863, 4776, -330, -3988, 
    -8517, -13038, -16824, -18909, -24933, -26269, -27205, -28571, -29911, 
    -31483, -31289, -27781, -27764, -24942, -24070, -20579, -15329, -13307, 
    -8270, -4467, -1055, 5290, 7234, 12779, 17150, 21679, 22834, 25626, 
    29385, 30918, 30325, 31233, 29606, 29505, 29301, 25182, 24656, 21159, 
    17059, 13370, 8865, 5625, 356, -4771, -8369, -12538, -17499, -21308, 
    -22890, -26049, -29235, -29071, -29614, -29530, -30248, -29312, -26331, 
    -26196, -23306, -19800, -17243, -14764, -9225, -5805, -480, 4675, 7379, 
    12744, 15615, 19315, 22316, 25051, 27396, 31071, 30004, 31811, 30859, 
    30945, 28705, 25869, 23397, 20860, 16745, 14349, 10021, 4937, -1013, 
    -3445, -9371, -12887, -15890, -20572, -22884, -24620, -26903, -29269, 
    -31053, -32068, -29424, -30088, -28803, -25857, -23312, -21476, -18239, 
    -14634, -8955, -4436, 409, 4512, 9382, 11301, 14929, 19635, 22438, 24619, 
    26203, 27938, 30155, 30853, 30063, 30098, 29923, 26302, 23436, 21499, 
    17212, 13343, 9117, 5391, 305, -3640, -8667, -10917, -15503, -19807, 
    -22194, -24928, -27275, -30336, -30598, -30962, -30379, -31338, -29110, 
    -25890, -24208, -20604, -17508, -14578, -9707, -3766, -321, 2680, 7741, 
    11660, 15336, 19749, 23503, 24383, 27820, 29731, 30884, 29598, 31087, 
    31416, 27363, 27875, 25218, 21040, 17682, 13320, 10057, 5957, 1867, 
    -2805, -7078, -12286, -16733, -20318, -22408, -24924, -26431, -28747, 
    -30036, -30820, -31844, -31058, -30133, -28140, -24143, -20645, -17495, 
    -13483, -9214, -6444, -2661, 3929, 7398, 10973, 14034, 19512, 22274, 
    24648, 27684, 27222, 29838, 29502, 29131, 30395, 29107, 27821, 25738, 
    22333, 17554, 14039, 10237, 6337, 2970, -1123, -7689, -11008, -15199, 
    -18403, -21682, -25736, -28690, -28117, -30291, -31441, -29024, -31490, 
    -29171, -26009, -25893, -21050, -18598, -14190, -10705, -5291, -804, 
    2002, 6453, 9873, 15340, 17704, 22380, 24327, 27234, 29293, 29209, 31118, 
    31592, 30172, 27482, 26333, 24320, 21033, 18557, 13834, 10716, 7046, 
    3404, -1200, -7164, -10254, -14194, -18123, -21110, -24803, -27467, 
    -28190, -29531, -30153, -30897, -31507, -29165, -25757, -24521, -22782, 
    -18251, -15172, -10069, -5833, -1173, 2047, 7526, 9894, 13148, 17456, 
    20904, 24673, 26588, 28014, 30583, 32452, 29816, 30430, 29372, 27364, 
    24032, 22190, 18625, 14783, 10319, 7051, 3642, -2385, -5006, -8691, 
    -14271, -19344, -21857, -23078, -25482, -29874, -31473, -30491, -31338, 
    -29209, -29019, -27467, -24667, -22642, -18244, -14324, -12674, -8474, 
    -4003, 1743, 5331, 10380, 13714, 17568, 19760, 22787, 26431, 27403, 
    29301, 30754, 30649, 29416, 27759, 27291, 24840, 21399, 20840, 15747, 
    10950, 8715, 2614, -1440, -5550, -10590, -13052, -17889, -20824, -23012, 
    -26311, -27129, -30849, -29970, -31290, -30835, -29970, -27896, -25293, 
    -23644, -18958, -15223, -11788, -6733, -4840, 1100, 6794, 8803, 15221, 
    16977, 21039, 24092, 25545, 28913, 29730, 29633, 31124, 29357, 29123, 
    28348, 24044, 22344, 20510, 14624, 12688, 8632, 4692, -1445, -4900, 
    -11190, -13295, -17865, -20413, -23133, -26395, -26590, -28520, -29732, 
    -30294, -29072, -30768, -27685, -26288, -22547, -19866, -16351, -12177, 
    -7323, -4313, 106, 5975, 8373, 14033, 16759, 19896, 23212, 25621, 28111, 
    28936, 30140, 31533, 29736, 27892, 26311, 25957, 22796, 20918, 15963, 
    12282, 7428, 4844, 179, -5536, -9722, -11995, -15297, -21290, -22833, 
    -27015, -28768, -29570, -29117, -30179, -30423, -29188, -29336, -25832, 
    -23146, -18643, -16365, -11458, -9912, -2819, -232, 3227, 7664, 12427, 
    15843, 18373, 23242, 25864, 28357, 29020, 31101, 30521, 29804, 30925, 
    28805, 25817, 23427, 21370, 16702, 14757, 9346, 4368, -151, -2283, -9356, 
    -13315, -17256, -19509, -23740, -27273, -27258, -28299, -30460, -31477, 
    -30596, -29836, -27902, -26045, -24772, -20417, -17914, -13024, -8753, 
    -5456, -1211, 4417, 9201, 12240, 15944, 19274, 21486, 24906, 28737, 
    29557, 30872, 31354, 30590, 29056, 28396, 26269, 22553, 20308, 16691, 
    13461, 9692, 4779, 766, -3722, -7875, -12836, -14811, -19682, -23824, 
    -27303, -27851, -28663, -30734, -30290, -31203, -31086, -27437, -25484, 
    -24892, -22277, -18324, -12221, -10340, -5996, -523, 4110, 8106, 11896, 
    16283, 19554, 21933, 26084, 28996, 29239, 30596, 30221, 30603, 28372, 
    27703, 26142, 23968, 19879, 17069, 14309, 10945, 5086, 2061, -3578, 
    -8301, -11459, -14775, -19468, -21683, -26123, -27313, -28298, -31214, 
    -31226, -31643, -29989, -28773, -25762, -24131, -19627, -18272, -14155, 
    -8791, -4456, -2382, 1329, 7491, 10738, 13679, 18784, 23901, 24785, 
    28154, 28994, 31103, 31244, 30784, 30507, 27084, 26219, 24890, 20301, 
    18158, 14845, 11167, 6363, 1049, -3113, -6658, -10332, -15586, -19829, 
    -23274, -23887, -27658, -28276, -30098, -29705, -31233, -29587, -29438, 
    -26973, -24017, -20827, -19286, -15007, -10316, -5667, -2877, 3142, 6135, 
    10938, 15741, 19347, 21881, 24407, 26527, 28773, 29354, 31858, 29210, 
    29904, 29318, 26800, 24767, 21527, 18793, 15847, 9433, 6117, 2790, -2919, 
    -7460, -12126, -14758, -18272, -21920, -24576, -27559, -29752, -29240, 
    -29738, -29854, -31209, -27963, -27491, -25195, -21458, -17822, -14969, 
    -11515, -6692, -1061, 565, 5123, 11111, 14686, 18366, 22375, 24680, 
    27254, 29706, 29923, 31026, 30915, 30064, 30218, 26636, 25851, 20515, 
    19096, 14984, 10757, 7722, 1943, -1003, -6617, -11112, -14878, -18127, 
    -21547, -23673, -27869, -29145, -29695, -31098, -31034, -31100, -30596, 
    -28147, -24198, -21883, -19297, -14159, -11209, -8052, -2777, 2301, 6220, 
    9202, 13203, 16668, 21367, 25003, 27647, 27970, 30757, 31138, 31909, 
    30129, 28170, 27299, 25493, 21634, 18824, 15504, 11104, 7975, 2999, 
    -3046, -5942, -9001, -14541, -16927, -21553, -25451, -25939, -29374, 
    -29708, -32530, -29967, -29213, -27427, -27177, -26251, -21940, -17596, 
    -14844, -11084, -7928, -3564, 1873, 5875, 10700, 12833, 17498, 22147, 
    23435, 27504, 27623, 29790, 29700, 29960, 30431, 29320, 29221, 23505, 
    23259, 19170, 15010, 13029, 7499, 3117, -2047, -4817, -9883, -13373, 
    -18603, -21592, -23822, -26010, -28221, -29007, -29593, -31169, -30715, 
    -29234, -27309, -25509, -21960, -19781, -16395, -12960, -8539, -3159, 
    679, 4287, 9150, 13578, 17019, 19598, 24906, 25307, 27686, 31106, 31927, 
    30976, 29764, 28941, 27289, 25166, 23310, 20147, 17092, 11641, 7059, 
    3614, -1202, -5934, -9836, -13673, -17014, -21002, -22559, -24792, 
    -26651, -29696, -30522, -31649, -30490, -29026, -27793, -24660, -22318, 
    -20737, -16537, -12624, -7426, -3003, 1375, 4262, 8947, 13004, 17620, 
    20899, 23678, 25592, 28170, 31169, 29804, 29651, 29960, 29239, 27314, 
    26212, 22364, 19467, 17169, 11224, 7271, 5420, -332, -6009, -8375, 
    -12779, -16880, -20688, -22932, -26696, -27885, -29867, -29768, -29807, 
    -31152, -28212, -28577, -25868, -23499, -21096, -16988, -11667, -8685, 
    -4203, 791, 3759, 8773, 12622, 17421, 21093, 22258, 26378, 27833, 27878, 
    31188, 30433, 32206, 29477, 27045, 26537, 24344, 20615, 17037, 12162, 
    9761, 4063, -325, -4435, -8755, -13454, -16334, -19631, -23533, -26506, 
    -27241, -29353, -30650, -30962, -30462, -30183, -29131, -26074, -22716, 
    -22284, -15975, -14253, -9401, -6017, -2102, 3503, 7861, 14094, 16799, 
    20880, 22593, 25576, 27314, 29150, 30134, 31081, 30912, 29197, 27768, 
    25887, 23101, 19091, 17528, 14936, 10095, 5529, 1704, -2724, -7074, 
    -11423, -15235, -19679, -22489, -25587, -27719, -30135, -31554, -30016, 
    -30611, -28604, -27778, -26395, -22726, -20130, -18721, -14639, -9901, 
    -6734, -657, 4375, 7904, 11032, 16621, 18677, 22639, 26882, 27855, 27982, 
    31134, 30990, 30438, 29041, 29906, 26857, 23519, 21191, 18467, 13861, 
    9615, 4714, 1172, -2487, -7149, -12543, -16181, -19152, -22137, -25240, 
    -26940, -29472, -32047, -31542, -30482, -31133, -29257, -26468, -23595, 
    -20347, -17328, -12429, -10886, -5065, -2682, 4350, 6680, 11433, 16034, 
    19687, 22128, 25772, 27617, 29478, 30122, 31286, 30228, 29108, 28101, 
    27659, 25179, 19538, 18138, 13687, 11281, 6159, 1536, -1970, -6696, 
    -11578, -14351, -18592, -20557, -24453, -27875, -29047, -29766, -29553, 
    -30071, -29218, -27529, -27036, -22765, -21450, -17793, -14652, -11032, 
    -5903, -2571, 2682, 6766, 11043, 13622, 19214, 22054, 24145, 27222, 
    30767, 29988, 30513, 30829, 30746, 29151, 26120, 24991, 22564, 18097, 
    12674, 11110, 5406, 2105, -2758, -7357, -10365, -15038, -19242, -21104, 
    -25884, -26745, -29067, -31395, -30496, -29565, -28640, -29865, -27202, 
    -25279, -21467, -18910, -15066, -10950, -5163, -2467, 1687, 6248, 10894, 
    13923, 18524, 21699, 25062, 27034, 27646, 30312, 29579, 29729, 30059, 
    28647, 27012, 25168, 21295, 19730, 16268, 10530, 6826, 899, -1457, -7684, 
    -9220, -14760, -18098, -21014, -24863, -26673, -28667, -29149, -32047, 
    -30845, -29991, -30903, -28010, -25385, -21283, -18885, -14713, -11744, 
    -8196, -2850, 279, 6456, 9151, 15963, 18853, 21023, 25045, 27850, 30434, 
    30249, 30364, 30289, 30378, 29866, 27575, 25158, 23683, 20315, 15312, 
    10740, 5942, 2882, -1266, -6350, -10516, -13916, -17075, -21923, -24133, 
    -26541, -28763, -28269, -31535, -31692, -31040, -29944, -26758, -25514, 
    -22612, -18528, -15782, -12163, -7831, -3296, 570, 5602, 9914, 14914, 
    16859, 20620, 23386, 27197, 26892, 28964, 29974, 30773, 28974, 29158, 
    27779, 24762, 22378, 18325, 14307, 12428, 8224, 4349, -741, -3900, -9121, 
    -14422, -17091, -21391, -23809, -25921, -27580, -30304, -30962, -30217, 
    -29560, -29290, -27392, -24677, -22577, -19124, -15932, -12045, -7632, 
    -3747, 2385, 5539, 8246, 12979, 19045, 21188, 25133, 26829, 30142, 29464, 
    30040, 32313, 30492, 28044, 28474, 26761, 24189, 20180, 16422, 13041, 
    8514, 4068, -506, -4968, -10555, -13917, -18485, -20479, -23496, -26546, 
    -28378, -30485, -30869, -29759, -30550, -29194, -28024, -24818, -22379, 
    -18822, -16733, -12343, -8690, -4314, 1144, 4418, 9670, 12305, 16794, 
    20551, 22223, 26114, 28955, 30311, 30003, 30855, 30754, 29284, 29019, 
    27385, 22712, 21258, 17739, 11377, 8827, 4196, -761, -5460, -8797, 
    -12128, -18020, -20166, -22933, -26558, -28172, -31130, -30488, -30672, 
    -30609, -29122, -28398, -26006, -24795, -19253, -15079, -11797, -8585, 
    -5553, 813, 4427, 8389, 13226, 15370, 19954, 24651, 24665, 26932, 28474, 
    31554, 31920, 29224, 28574, 28343, 25759, 22952, 19451, 16563, 13586, 
    10421, 2958, 748, -3535, -7352, -11880, -16099, -20163, -23142, -26842, 
    -26426, -30278, -30344, -30370, -30000, -29485, -28103, -25992, -24377, 
    -20953, -16475, -11823, -8604, -3431, -839, 5426, 7770, 12047, 17716, 
    20118, 23135, 26428, 28732, 29497, 30932, 29922, 29329, 31012, 29387, 
    27002, 22672, 22412, 18355, 13463, 9251, 4311, 2487, -3273, -7748, 
    -12834, -16690, -20178, -22216, -26228, -28368, -28290, -29509, -31636, 
    -29666, -30002, -29176, -26088, -23426, -21218, -17715, -14126, -9764, 
    -6106, -269, 3922, 9239, 11916, 15525, 18767, 21258, 25779, 27768, 28021, 
    32135, 31677, 30509, 30170, 29460, 27368, 24394, 19314, 16861, 13060, 
    8435, 3806, 2119, -3327, -6313, -11534, -14125, -19726, -23256, -24932, 
    -27419, -29106, -31106, -30028, -30670, -30467, -29471, -25867, -23147, 
    -20230, -17242, -12987, -9342, -4604, -1914, 3242, 6528, 9910, 14846, 
    19320, 22426, 26193, 28377, 30565, 30460, 30857, 29526, 31364, 29561, 
    26106, 25503, 22122, 17510, 15572, 10806, 5070, 954, -3516, -6968, 
    -11643, -15386, -18403, -23374, -24607, -26986, -28388, -30831, -30933, 
    -30222, -30058, -30104, -28063, -23111, -21830, -18252, -15208, -11490, 
    -6129, -1358, 1811, 6647, 10843, 14525, 17749, 22169, 25378, 28652, 
    29245, 30564, 32476, 30956, 31690, 29574, 27109, 23426, 22784, 19505, 
    13888, 10956, 6630, 145, -4142, -7302, -9427, -16205, -18623, -22599, 
    -24980, -27759, -29364, -29245, -32125, -31818, -29099, -27851, -28414, 
    -25045, -23115, -18633, -15884, -11123, -5695, -2031, 2343, 7608, 11412, 
    13331, 18053, 21339, 25185, 28052, 29430, 29046, 32195, 30054, 28724, 
    28851, 28427, 24216, 21845, 18826, 15569, 10148, 7716, 2210, -1907, 
    -6517, -10795, -14609, -17143, -21610, -24874, -27137, -29985, -30987, 
    -30125, -30581, -29335, -29407, -27384, -23546, -22012, -18926, -15445, 
    -11334, -6816, -3218, 1119, 6758, 11099, 14645, 18145, 21321, 25497, 
    26751, 28316, 29586, 32072, 30048, 28736, 28216, 28782, 25368, 23555, 
    18501, 14862, 11278, 7707, 2377, -1865, -6083, -9975, -15203, -18480, 
    -21916, -23714, -26932, -28085, -28899, -30934, -30193, -28880, -29199, 
    -26776, -24446, -23409, -19073, -15809, -12140, -7704, -4111, 2009, 4744, 
    8963, 13175, 18540, 20714, 23443, 26435, 27992, 30391, 30552, 29836, 
    29153, 29563, 27760, 25384, 22695, 18968, 14755, 11426, 7080, 2740, -700, 
    -5038, -9472, -14527, -17704, -20662, -23508, -26009, -28949, -31402, 
    -30154, -31152, -31254, -28506, -28839, -24832, -22422, -19574, -17037, 
    -11389, -9337, -2525, 895, 5104, 9667, 14228, 18915, 19293, 23820, 26737, 
    28601, 28633, 31407, 30628, 29689, 29129, 29415, 26995, 22025, 19602, 
    17474, 11403, 7830, 4557, 351, -3565, -7493, -14102, -16764, -19556, 
    -23554, -25061, -28112, -28171, -30535, -29252, -29637, -29792, -28032, 
    -24622, -23157, -19210, -16408, -11964, -8449, -3812, 685, 5598, 9583, 
    13619, 16112, 19536, 23711, 27017, 28776, 30262, 30822, 30424, 31324, 
    29714, 27880, 26312, 23983, 19777, 16396, 11218, 7613, 3964, -421, -5094, 
    -9146, -12563, -17971, -20659, -23399, -26056, -27681, -30139, -30837, 
    -30068, -30475, -29592, -28573, -25039, -22963, -19102, -15732, -11978, 
    -8520, -4984, 577, 4593, 7681, 12072, 15272, 19906, 23887, 25704, 27538, 
    28190, 31193, 29681, 30922, 29098, 27505, 26747, 23835, 19414, 16677, 
    12815, 8913, 4682, -1598, -3366, -9024, -11919, -16026, -18774, -22397, 
    -26323, -27883, -28368, -30737, -30918, -30935, -29355, -27466, -25610, 
    -22435, -21427, -15599, -12988, -9851, -4612, -1566, 3098, 8158, 13615, 
    15223, 19298, 22184, 24992, 27649, 30577, 31122, 30662, 30895, 31293, 
    29429, 27184, 23714, 21000, 16486, 12626, 8322, 4966, 605, -2980, -9195, 
    -10661, -15800, -19590, -23649, -24794, -28808, -29191, -30392, -30491, 
    -29888, -29305, -29140, -25559, -24246, -20828, -17817, -15029, -9863, 
    -5408, -1478, 2387, 8970, 11790, 16671, 19053, 21969, 25327, 28775, 
    28336, 30471, 30464, 30901, 30094, 29358, 27160, 24808, 21425, 18865, 
    15009, 10576, 5462, 1338, -3551, -8591, -10986, -15627, -19451, -22860, 
    -24845, -26799, -29610, -30476, -31204, -29644, -28609, -27500, -27606, 
    -24695, -19648, -16744, -14132, -9684, -5652, -677, 3129, 7379, 12328, 
    16347, 20608, 22616, 25237, 25970, 28250, 31050, 31055, 30716, 31024, 
    28452, 27659, 22941, 22712, 17848, 14100, 11027, 6852, 932, -1813, -6428, 
    -10933, -14378, -18632, -21032, -24019, -26909, -28150, -30780, -30387, 
    -30418, -29909, -29308, -26727, -23219, -22275, -18260, -13891, -9604, 
    -6656, -1665, 3988, 6945, 10641, 14237, 18774, 23108, 26514, 27128, 
    29240, 29032, 29391, 30665, 30035, 30119, 25621, 25044, 22893, 17099, 
    14049, 10648, 7013, 725, -1986, -6151, -10637, -15160, -19571, -22069, 
    -23662, -26654, -28420, -31216, -31375, -29164, -28809, -29443, -26590, 
    -24627, -22169, -18444, -14226, -10799, -5140, -3589, 1703, 6555, 11558, 
    14513, 17838, 21259, 25300, 27181, 29251, 30223, 32310, 29648, 30576, 
    28554, 27356, 26277, 21901, 18958, 15745, 11141, 7410, 2281, -1368, 
    -6249, -11270, -13947, -17791, -21165, -25449, -27480, -27624, -31391, 
    -29828, -30544, -31039, -29406, -27339, -24329, -22459, -19656, -16158, 
    -11741, -7503, -2299, 405, 6450, 9737, 14310, 18043, 22166, 24064, 26531, 
    27748, 29849, 30130, 32366, 31054, 27878, 28475, 23578, 21159, 18791, 
    16643, 11474, 7344, 2248, -1674, -5155, -10609, -13945, -16665, -20888, 
    -24511, -27282, -28883, -30634, -29701, -31186, -31246, -29113, -27450, 
    -25149, -22010, -19884, -15421, -10917, -7634, -4474, 988, 4046, 8444, 
    15343, 19052, 20929, 23663, 25642, 29682, 28777, 30003, 30827, 31217, 
    29712, 26345, 24862, 22694, 20254, 15938, 11741, 9370, 4215, -1441, 
    -4693, -10705, -13266, -17351, -20531, -24406, -27006, -28747, -28549, 
    -30509, -31631, -31144, -28880, -28044, -25451, -21415, -20089, -15982, 
    -11982, -7975, -3372, 1684, 4825, 8691, 13654, 19068, 21795, 22692, 
    25004, 29539, 29841, 30483, 31984, 30279, 29972, 28183, 24680, 23854, 
    20923, 17319, 12620, 6739, 2872, -552, -6238, -10554, -12494, -17048, 
    -21503, -23458, -26067, -28567, -29902, -30686, -29343, -30929, -29957, 
    -27941, -25275, -23656, -18406, -16864, -11879, -8020, -3671, 74, 3579, 
    9567, 14153, 17330, 19873, 24116, 26544, 29863, 29774, 30595, 30490, 
    30408, 28776, 27568, 26022, 23225, 20740, 15682, 12414, 9232, 4620, 553, 
    -5421, -8906, -13028, -17394, -21543, -24867, -26069, -28800, -30586, 
    -29421, -29675, -30905, -29713, -26987, -27101, -23580, -20409, -16906, 
    -12813, -8864, -4002, -1482, 5991, 8053, 13551, 16131, 21278, 23926, 
    26775, 28228, 30086, 30638, 31480, 31946, 28218, 27119, 24752, 24111, 
    20270, 18340, 13322, 8239, 4923, -731, -2853, -9557, -12028, -17846, 
    -19147, -22069, -25229, -27744, -29325, -30977, -32077, -31652, -28968, 
    -27924, -27398, -23124, -20681, -16168, -13301, -10448, -5273, -643, 
    3078, 8107, 11996, 16530, 19989, 22634, 26960, 28967, 29987, 30556, 
    32064, 30072, 29653, 27622, 26538, 23902, 20415, 17160, 13614, 7464, 
    4070, 362, -3694, -7647, -11456, -17303, -20399, -23437, -26943, -26558, 
    -30143, -30027, -30374, -30796, -30094, -29025, -26134, -23717, -19869, 
    -17776, -13307, -11242, -5835, -343, 3449, 7845, 10570, 17445, 18945, 
    22688, 25286, 29171, 30462, 31719, 31492, 30429, 30488, 28359, 26419, 
    24376, 19697, 18525, 12949, 10349, 6871, 1722, -4089, -7586, -12043, 
    -16216, -19114, -23048, -23555, -26981, -27845, -30535, -31042, -29965, 
    -29786, -28877, -25138, -23030, -20843, -18629, -14059, -10359, -4953, 
    -941, 2911, 7651, 12247, 16221, 19555, 21479, 24111, 27484, 28158, 30443, 
    31100, 31234, 30210, 28887, 26728, 23993, 20762, 18387, 15218, 10935, 
    6335, 990, -1423, -6434, -11625, -15294, -20192, -22477, -25308, -25695, 
    -28944, -30125, -29196, -30599, -29774, -29704, -24968, -25854, -21458, 
    -18074, -12503, -10148, -6724, -2585, 4080, 6110, 10651, 16479, 18493, 
    21398, 25055, 28581, 28205, 30441, 31839, 32084, 30102, 28375, 25395, 
    25246, 20873, 17636, 15398, 11413, 5742, 1711, -3107, -6963, -9824, 
    -14703, -18782, -21967, -23707, -26622, -30335, -30216, -29774, -32164, 
    -30571, -29521, -28132, -24323, -21392, -17321, -13733, -11498, -7002, 
    -2203, 2502, 7136, 9447, 14104, 17607, 21892, 23620, 25730, 29362, 29559, 
    31313, 30640, 30516, 28367, 27063, 24071, 21335, 19524, 15048, 12019, 
    7174, 3449, -2815, -5902, -11232, -15692, -18776, -21824, -25332, -26524, 
    -27597, -31074, -32274, -30866, -29568, -28372, -27216, -23367, -23655, 
    -17450, -14767, -9645, -8028, -2684, 1426, 5226, 10162, 15780, 17810, 
    22685, 24675, 25666, 28097, 29309, 31995, 32420, 31571, 29193, 28480, 
    25937, 22825, 20735, 14012, 12053, 7336, 3083, 32, -6031, -9680, -14919, 
    -18780, -22331, -25891, -26334, -29620, -29327, -31538, -30502, -31283, 
    -27283, -26557, -25807, -22975, -17859, -14063, -11814, -6323, -3060, 
    815, 5212, 9207, 14288, 18299, 20707, 24452, 26299, 28017, 28392, 29516, 
    30947, 31395, 29827, 26701, 24552, 24147, 19486, 17159, 12409, 6508, 
    3377, -2205, -5390, -7956, -14837, -17983, -20271, -23623, -25507, 
    -29000, -29528, -30658, -30483, -30883, -29639, -27471, -23771, -21875, 
    -19113, -15694, -12621, -6342, -2815, -499, 4615, 9992, 13848, 17240, 
    22082, 23121, 25065, 27422, 29334, 31575, 32126, 31668, 29153, 28765, 
    24774, 24357, 19243, 17347, 11749, 9216, 3584, -1144, -6455, -8857, 
    -13163, -16686, -21488, -23486, -26544, -29312, -29037, -31078, -31835, 
    -31242, -29458, -27567, -25594, -21971, -18491, -16523, -12693, -7400, 
    -4727, -1228, 4630, 9268, 12219, 17794, 20558, 23289, 26766, 27786, 
    29087, 29712, 29544, 31021, 28734, 27848, 26169, 24431, 20300, 16749, 
    11936, 8897, 3170, 862, -4393, -8684, -12275, -17323, -20890, -24305, 
    -24486, -28129, -28620, -30923, -30074, -31328, -29286, -26384, -24887, 
    -23537, -19628, -15230, -14468, -10513, -4578, -331, 5122, 10202, 13398, 
    16174, 20198, 24131, 25669, 28094, 30517, 30833, 31743, 29607, 29229, 
    27503, 25513, 22595, 20576, 18551, 13233, 8969, 3099, 388, -3018, -8701, 
    -11609, -16242, -19861, -21997, -24074, -27776, -29953, -29675, -31892, 
    -30608, -29422, -27616, -26451, -23600, -21268, -16012, -12646, -10194, 
    -4697, -242, 4937, 7755, 10710, 16409, 18685, 24730, 24056, 26525, 30102, 
    31914, 30718, 31236, 30239, 28497, 26587, 22784, 21774, 16210, 12941, 
    8473, 4703, 191, -4029, -7646, -12196, -15423, -18901, -22966, -26321, 
    -27104, -29702, -31363, -31519, -30076, -31265, -28228, -26040, -22311, 
    -20096, -17190, -14265, -8098, -4637, -816, 3668, 6618, 12127, 15488, 
    19301, 23081, 26939, 27436, 30389, 31127, 32126, 29486, 29634, 28766, 
    28109, 23183, 21428, 17232, 13238, 10513, 4159, 398, -2559, -6406, 
    -11978, -15221, -18519, -21076, -25261, -27367, -29671, -30769, -30325, 
    -29872, -31390, -29437, -27537, -23952, -19896, -17843, -12652, -11610, 
    -5967, 363, 2969, 7556, 10718, 17155, 21043, 22343, 24656, 26496, 30598, 
    28757, 30570, 32201, 30215, 28719, 26715, 23714, 21976, 17841, 12997, 
    10810, 5930, 2851, -2652, -7314, -11305, -15392, -18671, -23683, -24664, 
    -26929, -29908, -31214, -29691, -29314, -29735, -28744, -27565, -24843, 
    -21769, -19044, -14287, -9596, -5883, -2492, 1507, 6879, 10966, 16077, 
    17974, 21085, 25500, 26441, 28394, 29596, 31060, 31057, 30293, 28266, 
    27253, 23302, 21846, 18004, 14663, 10999, 6571, 3281, -2119, -6194, 
    -11174, -14650, -18690, -21811, -24086, -26162, -28147, -31714, -30219, 
    -29386, -30505, -29925, -25866, -25044, -20635, -19784, -15668, -10836, 
    -6835, -1326, 1119, 7088, 11826, 14557, 17513, 20529, 25662, 27056, 
    28957, 29288, 31115, 30940, 29365, 29217, 27295, 24465, 21608, 18485, 
    15098, 12036, 7188, 2441, -3154, -6241, -11925, -14602, -17683, -21032, 
    -22938, -27008, -27504, -30189, -31399, -31808, -29942, -28273, -28376, 
    -24998, -21693, -19211, -15623, -11029, -7237, -1249, 2767, 7591, 10697, 
    13511, 17437, 21584, 23410, 26359, 28300, 29350, 31519, 32146, 31341, 
    29389, 26464, 23785, 21852, 19311, 15380, 10991, 7929, 1197, -2058, 
    -5210, -10510, -12499, -17386, -20404, -25018, -27194, -29124, -31042, 
    -29845, -30819, -29853, -29342, -27475, -24617, -22364, -19332, -14492, 
    -10808, -6236, -3324, 1981, 6608, 8840, 12649, 17374, 21403, 24980, 
    27106, 29120, 30317, 29118, 29611, 29806, 29866, 29404, 25220, 22548, 
    19758, 14551, 10967, 5866, 4861, -812, -4427, -9866, -13923, -17706, 
    -20987, -24110, -26598, -29177, -29904, -29648, -30714, -32193, -29314, 
    -27420, -26707, -21930, -18519, -17711, -12885, -7053, -3409, -603, 4527, 
    10481, 14081, 16201, 21115, 24751, 25320, 28988, 30242, 30486, 31090, 
    29715, 28136, 26919, 25736, 23849, 19736, 16510, 11083, 7966, 3702, 266, 
    -6661, -9395, -12904, -16645, -21299, -23089, -26312, -28019, -29945, 
    -29937, -30828, -30240, -28899, -27506, -25373, -23888, -19065, -16532, 
    -11882, -9110, -3133, 1064, 4823, 9769, 11833, 18690, 21396, 23763, 
    25569, 29399, 28547, 30158, 32085, 29731, 30202, 27147, 25696, 22510, 
    20738, 16952, 13488, 8550, 5460, -294, -4751, -9473, -13356, -16542, 
    -20991, -24382, -26272, -28169, -29537, -30357, -30448, -29419, -28276, 
    -27092, -25974, -23244, -19714, -15890, -13812, -8460, -3852, -1145, 
    2842, 8345, 13893, 16379, 19523, 22519, 26565, 26868, 31302, 31095, 
    29164, 29357, 31099, 27933, 27123, 23403, 20436, 17066, 12372, 9060, 
    3234, -689, -5705, -8731, -12093, -17197, -19198, -22840, -27236, -26953, 
    -29832, -31270, -30306, -31663, -28339, -27219, -26711, -23439, -22264, 
    -16112, -13297, -10339, -5028, 890, 3252, 7156, 11327, 14630, 19514, 
    22997, 25759, 26850, 28845, 31647, 30846, 29728, 29906, 29543, 25635, 
    25240, 20413, 17284, 13604, 10118, 5075, 373, -2795, -7597, -11538, 
    -15305, -19198, -24371, -25489, -27111, -29213, -30492, -32626, -31959, 
    -30524, -28844, -25952, -24615, -21155, -18417, -14013, -9159, -6911, 
    -675, 3949, 7503, 11018, 16408, 18495, 22418, 25346, 28027, 29265, 29522, 
    31070, 30047, 30677, 27447, 27156, 23331, 21745, 18333, 15009, 8927, 
    4783, 1291, -4525, -8487, -11484, -14104, -19955, -22295, -25520, -28458, 
    -29900, -30283, -29999, -30881, -31254, -27660, -26183, -24023, -20772, 
    -17317, -14644, -9828, -5987, -196, 2832, 5776, 11578, 15331, 17816, 
    22056, 26161, 27485, 29185, 31082, 30782, 31313, 29283, 27951, 25285, 
    23512, 22039, 17908, 13364, 11735, 6639, 582, -3822, -6720, -11099, 
    -16007, -17865, -22783, -24041, -25877, -29509, -31186, -31662, -32096, 
    -28538, -28831, -26739, -22753, -22137, -18764, -14760, -10654, -6443, 
    -2018, 4058, 7127, 11808, 15411, 18161, 21982, 24953, 27346, 28795, 
    31016, 29864, 31765, 28895, 28342, 26760, 24470, 21706, 18521, 12855, 
    8892, 6907, 1322, -2126, -7217, -11386, -13770, -18711, -22186, -25569, 
    -27206, -28602, -30257, -30023, -30634, -31019, -29191, -26785, -23222, 
    -21717, -17953, -13413, -10075, -6842, -3638, 2454, 5630, 10880, 15341, 
    19971, 21129, 24792, 27313, 28886, 30405, 30249, 31593, 29756, 29611, 
    25893, 24885, 21972, 19322, 15561, 11608, 5932, 1503, -937, -4739, 
    -10386, -15221, -17046, -21770, -25472, -26937, -29049, -29484, -31791, 
    -30774, -30557, -29068, -26821, -25214, -22426, -18459, -15969, -11934, 
    -6733, -2686, 490, 6708, 10011, 15630, 19527, 20770, 25544, 26461, 27404, 
    29007, 30778, 31297, 30099, 29218, 27130, 24217, 22400, 19083, 15333, 
    10484, 6138, 3348, -1616, -5448, -10503, -14005, -18846, -19638, -24593, 
    -25074, -28975, -29162, -31320, -31403, -29731, -30998, -26759, -26301, 
    -21749, -20723, -16190, -9845, -5972, -2417, 1406, 6313, 9729, 13550, 
    18125, 21691, 23582, 26442, 29121, 28742, 29333, 31530, 30472, 28965, 
    28239, 24975, 21816, 20654, 16455, 11307, 7627, 4632, 151, -6158, -10770, 
    -13330, -17979, -20603, -22973, -27080, -27887, -29508, -31032, -31280, 
    -29006, -29186, -28432, -24660, -23707, -18830, -15708, -12879, -8404, 
    -2177, -46, 4610, 8626, 13198, 17182, 20853, 24621, 26490, 29557, 30854, 
    30323, 30491, 31746, 28746, 28274, 24784, 22646, 19368, 14892, 12037, 
    7154, 3139, -1953, -5210, -9339, -15206, -15942, -21294, -23793, -26772, 
    -28450, -28896, -29346, -30906, -29945, -28650, -26866, -26301, -22123, 
    -21075, -16783, -13411, -8545, -3882, -166, 3619, 9374, 13660, 16720, 
    21187, 23023, 27607, 27564, 28694, 32261, 30578, 30708, 29534, 27293, 
    25434, 23078, 20137, 15977, 12367, 8284, 4506, 1046, -4088, -10311, 
    -14036, -16788, -21018, -24172, -26666, -28969, -28379, -30416, -30988, 
    -31111, -29819, -27349, -25558, -23272, -20503, -17488, -13771, -9860, 
    -5372, -426, 4380, 8729, 12232, 15331, 19527, 23363, 24626, 27712, 29179, 
    30371, 30915, 30697, 30063, 29480, 25925, 22380, 19050, 16631, 13061, 
    7743, 4322, 594, -3709, -7767, -12104, -16736, -19493, -23978, -25746, 
    -26135, -28966, -31074, -29451, -30310, -29188, -27970, -26868, -24302, 
    -20328, -17113, -14513, -8522, -5947, -739, 3629, 8413, 13023, 15477, 
    19319, 24603, 26947, 28586, 29056, 30410, 31083, 30383, 28842, 28262, 
    24717, 23758, 21439, 18200, 12882, 10436, 6672, 1419, -5055, -7172, 
    -12203, -15634, -18961, -21486, -25235, -27930, -29328, -29613, -30591, 
    -31196, -30181, -29885, -26234, -23245, -20995, -16182, -12865, -8764, 
    -4561, -946, 3580, 8021, 11702, 14689, 19519, 23204, 24342, 28078, 29565, 
    30875, 30458, 29551, 29583, 29833, 27351, 23140, 20564, 17413, 12787, 
    8989, 5261, 1297, -4503, -6490, -10764, -15304, -19009, -23145, -25086, 
    -26221, -27942, -29238, -31396, -30915, -31176, -28603, -26218, -23662, 
    -21302, -18957, -13365, -9562, -6324, -2798, 1817, 7169, 10896, 15728, 
    18552, 21574, 26153, 28205, 29205, 30006, 30969, 30524, 30578, 27616, 
    26343, 24678, 22477, 16300, 13825, 9470, 4865, 1472, -1272, -6903, 
    -10884, -14482, -19648, -22735, -24915, -28155, -27604, -30337, -31670, 
    -29636, -31479, -29100, -28080, -24269, -21987, -16950, -13677, -11249, 
    -6150, -788, 2038, 7142, 11756, 14888, 17804, 22450, 26147, 25831, 29661, 
    30356, 29638, 29351, 29151, 28674, 27277, 24665, 21805, 18013, 14535, 
    9940, 5379, 2960, -3420, -6550, -10606, -15909, -17118, -21814, -25358, 
    -27769, -28810, -31010, -31049, -30843, -30061, -28370, -26371, -24543, 
    -21991, -17635, -14235, -10931, -5919, -2589, 2970, 6233, 10874, 15053, 
    18759, 20815, 25179, 26223, 27614, 29272, 32014, 29878, 29514, 29147, 
    25776, 24130, 23684, 18286, 15642, 11608, 6746, 2378, -1284, -6401, 
    -11093, -14480, -17644, -21508, -24113, -26694, -29428, -30033, -30374, 
    -30433, -30570, -27621, -27308, -25027, -21065, -19232, -14776, -12015, 
    -6877, -3364, 2336, 6265, 10321, 14979, 17761, 20639, 24213, 26980, 
    29388, 30270, 32095, 30068, 28748, 29984, 26795, 25384, 22458, 19712, 
    14542, 11968, 7580, 2829, -1666, -6902, -9754, -15014, -18672, -22553, 
    -24134, -26174, -28761, -30296, -31628, -31595, -29351, -27459, -28781, 
    -24214, -20906, -19009, -15226, -12838, -6401, -3276, 2252, 5000, 9707, 
    13611, 17714, 21935, 24663, 26721, 28194, 28650, 30614, 31219, 29508, 
    28887, 26460, 24199, 22653, 20291, 16799, 11074, 7184, 2918, -2243, 
    -7043, -9395, -13598, -17756, -19998, -24795, -25428, -30128, -31092, 
    -30550, -30999, -31161, -29391, -28054, -25631, -22900, -20133, -17086, 
    -13266, -8856, -2218, 583, 5587, 9412, 13922, 17992, 20981, 24323, 25538, 
    27531, 29670, 31474, 31086, 30874, 29261, 28424, 26779, 22531, 18957, 
    16057, 11491, 9024, 4736, 485, -5871, -8434, -12458, -16161, -21708, 
    -23280, -26286, -28421, -30574, -29219, -30753, -30395, -28098, -28007, 
    -25994, -22443, -19565, -15580, -12073, -7785, -2761, -732, 4106, 7509, 
    12676, 17400, 21660, 24486, 26879, 29110, 29322, 29927, 30179, 30361, 
    29220, 26696, 25406, 22420, 20652, 16214, 11943, 8178, 3836, 838, -4470, 
    -9073, -11973, -17053, -20728, -24223, -26704, -29200, -30668, -31582, 
    -31399, -31649, -29462, -26365, -25198, -23215, -19771, -17552, -12567, 
    -7446, -3877, 508, 3871, 9795, 13001, 16695, 21117, 22990, 27315, 28068, 
    29574, 29399, 31696, 31300, 29563, 26859, 26106, 24794, 19504, 16209, 
    12116, 7438, 4024, 292, -4555, -8489, -12920, -16454, -20583, -22627, 
    -26371, -27489, -28862, -31733, -31227, -31915, -28247, -28741, -25166, 
    -22763, -19533, -17119, -13174, -9873, -4887, -1420, 3964, 8246, 13181, 
    16722, 20131, 22297, 25230, 27144, 29829, 30644, 31285, 30262, 29619, 
    27911, 25265, 24145, 20409, 17616, 13101, 9623, 4435, 37, -3654, -7977, 
    -13356, -16040, -20261, -24194, -25075, -25931, -29901, -29859, -29972, 
    -32411, -30998, -27186, -25258, -23843, -20795, -18391, -14023, -8234, 
    -5973, -1619, 4764, 7578, 12429, 16045, 19444, 23500, 25152, 27033, 
    29558, 32062, 29628, 31235, 30326, 26968, 26601, 23585, 21248, 18171, 
    13463, 9380, 5550, 808, -2447, -9005, -11823, -15038, -19126, -21441, 
    -25401, -26187, -28839, -29258, -31045, -29513, -30816, -29749, -25979, 
    -24873, -22398, -17944, -14342, -9837, -5330, -1502, 3308, 6613, 12313, 
    15895, 17516, 21782, 26043, 27917, 30434, 31474, 30941, 32101, 31054, 
    27358, 26532, 25682, 21833, 18394, 14544, 9799, 6967, 277, -2863, -5825, 
    -11035, -16238, -18408, -22778, -24294, -26695, -29541, -29944, -30631, 
    -31436, -29256, -30279, -27313, -24468, -22064, -16866, -14184, -11027, 
    -6481, -939, 3672, 6369, 11838, 14894, 19481, 22774, 24662, 26628, 28264, 
    29352, 31260, 30031, 29789, 28724, 28234, 24759, 22644, 18030, 13601, 
    9345, 6640, 1648, -2783, -5827, -10399, -14970, -19321, -21822, -24510, 
    -26710, -28693, -30508, -30637, -30726, -29586, -27292, -27555, -24526, 
    -22758, -17770, -14727, -11446, -6671, -2565, 1629, 6011, 11782, 14961, 
    18379, 21490, 24258, 26924, 29719, 29632, 31527, 30341, 28678, 28331, 
    26033, 23990, 21145, 19771, 15924, 11683, 5436, 2300, -2892, -5643, 
    -10663, -15804, -17751, -21608, -23242, -26970, -29460, -28543, -30695, 
    -31610, -30511, -27791, -26526, -26022, -22048, -18418, -15161, -11287, 
    -7115, -2949, 1855, 6086, 10759, 15088, 16749, 21594, 23349, 25969, 
    29685, 30309, 30727, 29538, 31316, 29627, 26266, 26715, 23145, 18878, 
    15351, 9685, 5392, 3353, -2342, -6623, -9368, -12783, -16943, -22378, 
    -24568, -26931, -28410, -29296, -30415, -31236, -30100, -30178, -29240, 
    -25291, -21380, -19389, -13942, -10973, -8183, -3694, 1596, 5432, 10521, 
    14305, 16613, 21143, 23458, 27520, 28962, 31045, 30228, 30954, 29818, 
    28978, 26817, 25347, 22605, 19540, 17047, 11775, 7482, 3172, -750, -5525, 
    -10341, -12928, -19276, -21499, -25148, -26406, -28182, -29570, -30139, 
    -30509, -30212, -29036, -26782, -26328, -22236, -18695, -16376, -11323, 
    -7020, -3588, 1080, 5397, 11053, 12252, 18704, 21176, 22742, 27426, 
    28132, 28628, 29836, 30728, 30286, 29086, 27280, 24775, 21744, 19641, 
    17068, 11373, 6959, 2065, -669, -5127, -10403, -13552, -18546, -21641, 
    -21810, -27665, -27349, -29305, -30280, -31852, -29733, -30122, -26218, 
    -24455, -24721, -20408, -15464, -12263, -9247, -4856, -173, 5773, 9068, 
    13160, 17317, 20185, 22755, 25858, 28738, 29444, 31167, 30517, 31135, 
    28632, 26968, 24451, 23461, 20313, 16396, 12251, 9587, 4539, 1111, -5901, 
    -9844, -13131, -17986, -20027, -21553, -26383, -28210, -30045, -31099, 
    -29635, -29977, -30853, -26604, -27365, -22754, -20541, -16005, -12020, 
    -10059, -4310, 230, 4148, 7682, 13748, 16055, 19795, 23061, 25428, 28137, 
    30355, 30784, 32229, 30106, 28899, 28277, 25282, 23279, 21393, 17008, 
    12561, 8508, 3593, 396, -3981, -7864, -10972, -15730, -21460, -22886, 
    -26369, -27634, -30010, -31083, -30274, -30826, -30424, -28486, -26147, 
    -23055, -20533, -16428, -12638, -8847, -4481, -962, 4493, 8107, 14017, 
    15886, 20210, 23116, 24969, 27457, 30192, 30360, 32257, 30766, 30225, 
    27880, 26291, 24124, 22233, 17459, 13665, 9229, 5329, 1110, -5183, -8199, 
    -11279, -16035, -18817, -22925, -25657, -27773, -29346, -31566, -30043, 
    -31281, -28778, -28375, -27027, -23825, -19920, -16347, -14305, -10708, 
    -5746, -340, 3852, 8629, 11961, 14357, 19083, 23697, 26392, 27448, 29110, 
    30807, 30802, 31052, 29861, 26896, 26647, 23385, 20069, 17696, 14871, 
    9407, 4487, 1122, -4523, -7750, -12138, -15730, -20677, -23014, -24430, 
    -27854, -30072, -30250, -30307, -30466, -29921, -29237, -27249, -24979, 
    -21091, -18810, -12131, -8987, -6747, -1200, 1925, 7000, 11427, 14062, 
    17665, 21991, 25546, 27682, 29383, 31737, 30970, 30761, 29121, 28899, 
    27188, 24797, 19578, 17556, 15445, 9255, 6143, 978, -3149, -7078, -10540, 
    -14458, -17219, -21251, -25688, -26170, -28702, -30710, -29911, -31083, 
    -30180, -28139, -26405, -25291, -20971, -19416, -14768, -11082, -7232, 
    -2199, 4276, 8170, 11991, 15056, 18693, 21755, 23944, 27248, 29895, 
    30447, 29613, 30756, 30289, 27721, 27599, 24524, 20557, 18653, 16138, 
    9785, 6110, 442, -2427, -5832, -9849, -15690, -18545, -21030, -24718, 
    -28384, -28802, -31018, -31665, -31675, -30284, -29668, -26617, -23885, 
    -20650, -17273, -14944, -10309, -7486, -2007, 3712, 8185, 11933, 14577, 
    19901, 21605, 24474, 26892, 27924, 30138, 31018, 29789, 29154, 29762, 
    26951, 25949, 22619, 18034, 14421, 10592, 5836, 2337, -2416, -6436, 
    -10230, -14633, -19607, -20639, -24328, -27173, -28773, -30358, -31825, 
    -31054, -30427, -28722, -27350, -24173, -21915, -18710, -14895, -10720, 
    -6320, -2512, 1990, 4857, 8817, 15978, 16780, 20316, 24669, 26788, 28194, 
    30146, 30939, 32451, 30411, 29162, 25743, 24801, 21625, 18805, 14752, 
    11003, 5421, 2301, -2754, -4663, -9331, -13815, -18118, -20844, -25292, 
    -27041, -27605, -30281, -29487, -31255, -29703, -28770, -26554, -26618, 
    -22311, -18118, -15354, -11611, -7304, -2789, -87, 5963, 9277, 13869, 
    18432, 21641, 23096, 27699, 30092, 29299, 31258, 29461, 29499, 29134, 
    27419, 24907, 21181, 20871, 16992, 12725, 7842, 3313, -167, -5957, -9219, 
    -13903, -17389, -19342, -23117, -26883, -29167, -28672, -30640, -31267, 
    -29914, -29522, -28114, -23909, -22355, -20100, -14752, -11933, -8011, 
    -3278, 579, 5888, 9169, 13752, 16321, 19201, 25274, 25836, 27964, 28790, 
    30823, 29924, 28964, 27829, 27759, 26238, 22259, 18929, 17944, 12255, 
    7109, 2531, -36, -5314, -10262, -14724, -16050, -19308, -22789, -26341, 
    -27567, -29771, -31336, -30965, -30164, -28660, -28421, -25795, -23509, 
    -21305, -16668, -11306, -7215, -4624, 462, 6460, 8227, 12292, 16644, 
    21699, 23811, 26659, 26520, 28726, 29415, 30922, 29053, 30926, 29046, 
    26074, 24007, 19445, 16275, 14201, 9002, 4849, -1277, -4576, -9329, 
    -12874, -15745, -20937, -24848, -26832, -29895, -29376, -30478, -31646, 
    -29681, -29918, -26740, -26088, -22775, -21888, -16387, -11534, -8718, 
    -5027, 1398, 4276, 8681, 12085, 15882, 19355, 22795, 27094, 28502, 28081, 
    31223, 31317, 31440, 30683, 28494, 25528, 22125, 20187, 16984, 13010, 
    8540, 4875, 826, -3005, -10173, -13426, -17658, -21258, -21659, -25265, 
    -28956, -29737, -31452, -31206, -31148, -28285, -28283, -26521, -23291, 
    -21914, -17124, -12759, -8144, -5902, -1250, 4758, 9498, 12643, 16667, 
    19812, 22785, 26425, 27723, 30006, 30342, 31457, 30803, 29232, 27527, 
    25851, 24245, 20395, 17858, 13095, 9757, 3410, 1598, -1935, -7074, 
    -12972, -15633, -20234, -23352, -25752, -26994, -27668, -30638, -29543, 
    -30917, -30721, -28355, -26088, -24063, -20181, -17520, -13982, -9386, 
    -4372, -1762, 4594, 7926, 10570, 15937, 19429, 22852, 26970, 26879, 
    29136, 30777, 30463, 31157, 30253, 28963, 26197, 24012, 20729, 16838, 
    13478, 9959, 5942, 620, -2160, -7843, -12307, -16996, -19611, -22011, 
    -24590, -28807, -28465, -31649, -30536, -31074, -30687, -28062, -26462, 
    -23775, -21321, -19132, -14095, -8502, -5715, -720, 2893, 8302, 10947, 
    14032, 18774, 22097, 24570, 25716, 29536, 30959, 30797, 30653, 30197, 
    29800, 26740, 23269, 22735, 18909, 13339, 8815, 7039, 1336, -1779, -6781, 
    -10142, -15263, -20275, -22472, -24890, -27594, -29172, -29000, -30916, 
    -30611, -29808, -29135, -26184, -25085, -21991, -16868, -15319, -9178, 
    -7131, -2769, 4026, 7079, 11008, 15463, 18220, 22647, 23838, 26210, 
    29089, 29180, 32631, 29159, 30381, 29050, 27414, 24600, 22004, 19152, 
    15117, 9139, 5388, 2388, -2325, -6710, -10943, -15815, -18188, -21088, 
    -26406, -28189, -27620, -31099, -31008, -30711, -28935, -29240, -27038, 
    -23850, -22822, -19068, -13535, -9540, -5319, -1230, 605, 6497, 10537, 
    15653, 18855, 22451, 23794, 27536, 30650, 30457, 31613, 31515, 31116, 
    27350, 28106, 25333, 22214, 18384, 15487, 11402, 6656, 2050, -1761, 
    -6501, -11840, -15429, -18255, -21951, -23652, -26108, -28064, -29318, 
    -30396, -30766, -29402, -29429, -27294, -24129, -23368, -19510, -16307, 
    -10818, -6475, -2076, 630, 6401, 10124, 14366, 17104, 21169, 24360, 
    26403, 29345, 29613, 29756, 30830, 31172, 29931, 26431, 24662, 23422, 
    18850, 15269, 11594, 6429, 2209, -1567, -6601, -11436, -15297, -17632, 
    -22476, -23913, -27858, -27868, -29746, -29919, -32688, -30889, -28477, 
    -27089, -24493, -23367, -20388, -14745, -10957, -7643, -3687, 1686, 5289, 
    10881, 15047, 18280, 21719, 24632, 26582, 28572, 28838, 30286, 30189, 
    30651, 29714, 26666, 26390, 23477, 19451, 15255, 12259, 7672, 2111, -722, 
    -5292, -9347, -13196, -16686, -20849, -24945, -27073, -29928, -29061, 
    -32191, -30138, -29760, -29372, -28486, -24267, -22538, -18900, -16105, 
    -12325, -7692, -4309, -344, 4769, 9771, 13977, 16624, 19666, 24527, 
    26609, 28295, 29508, 32014, 30825, 31421, 28740, 26838, 23712, 22836, 
    18233, 15436, 11619, 8526, 3302, 128, -5195, -10156, -13614, -16864, 
    -22033, -22314, -25803, -26457, -29759, -30979, -29345, -31511, -28783, 
    -28222, -26366, -22810, -21486, -16627, -12381, -9047, -2226, 817, 3790, 
    10013, 14191, 17606, 21262, 24000, 24470, 28389, 31293, 30990, 31457, 
    31244, 30001, 28630, 26242, 23054, 20257, 17619, 11680, 9075, 4353, -159, 
    -4679, -8375, -13085, -17088, -18982, -23031, -27162, -27924, -28655, 
    -30166, -29593, -30636, -28414, -28448, -27022, -23280, -21652, -17611, 
    -12367, -8280, -4173, 423, 6012, 7685, 13646, 16984, 20211, 23750, 25692, 
    27636, 30758, 29443, 31052, 31028, 30706, 27388, 26334, 22860, 19682, 
    17864, 12225, 9831, 4829, 1336, -5318, -8919, -13242, -16479, -19049, 
    -22779, -24552, -28379, -29209, -32167, -29460, -31818, -29327, -26563, 
    -27368, -23402, -21032, -16728, -12857, -8529, -5115, -352, 5318, 6963, 
    12353, 16318, 20577, 21505, 25695, 28039, 29239, 30635, 31073, 31846, 
    28686, 26876, 27085, 23444, 20253, 17850, 14049, 7815, 4880, 157, -4285, 
    -7204, -11019, -17556, -20341, -22469, -24430, -29530, -29046, -30668, 
    -31610, -30781, -30655, -26933, -26067, -22800, -19837, -17273, -13663, 
    -9109, -5399, -1250, 3838, 7705, 11227, 14645, 18397, 21472, 24671, 
    27018, 30472, 29346, 29492, 29560, 30220, 28317, 27112, 23571, 20318, 
    18268, 13944, 9615, 6287, 1640, -2778, -8660, -12675, -16322, -17719, 
    -21967, -24846, -26464, -29369, -29133, -30555, -30612, -30761, -27807, 
    -27991, -25434, -21387, -18521, -14272, -9195, -7053, -539, 2345, 6125, 
    12408, 15260, 19733, 23826, 24511, 28525, 28039, 31012, 31793, 32273, 
    30215, 28633, 26215, 23893, 20672, 17567, 14723, 10947, 7183, 2674, 
    -3279, -7856, -11351, -16163, -18994, -22090, -25585, -26887, -29281, 
    -30665, -30081, -31356, -30768, -28168, -26160, -24836, -21601, -18186, 
    -14714, -12002, -4708, -2843, 3696, 6650, 11333, 14472, 19372, 21524, 
    25243, 26485, 29252, 29579, 30401, 30618, 28792, 29884, 26665, 24964, 
    20261, 17972, 13397, 10689, 6034, 2090, -1447, -7022, -11788, -15004, 
    -18868, -23189, -25158, -26144, -30337, -30258, -32002, -31774, -30873, 
    -27299, -26940, -22853, -20329, -19267, -15022, -10004, -8123, -2180, 
    2245, 8033, 11607, 15179, 17907, 21872, 24851, 26615, 28023, 29562, 
    32210, 31757, 31835, 28766, 26237, 24767, 21125, 19379, 14123, 10849, 
    7050, 2804, -1847, -5889, -10810, -16304, -18033, -22281, -24140, -27430, 
    -29896, -30882, -31209, -29618, -30982, -28709, -27123, -25570, -21519, 
    -17962, -15148, -11470, -6877, -2417, 1887, 6459, 12229, 14670, 16953, 
    20965, 24466, 26946, 27776, 30693, 31204, 30649, 31659, 28965, 26301, 
    25466, 21171, 18566, 15416, 12127, 7625, 3760, -1100, -5627, -9399, 
    -13295, -17530, -22323, -25090, -27493, -28595, -30900, -30671, -30183, 
    -29913, -28996, -26486, -26106, -22227, -19237, -15369, -11102, -7470, 
    -3211, 576, 5949, 9833, 13322, 17765, 20416, 23324, 27000, 28887, 29581, 
    31126, 29440, 29897, 29691, 27772, 24136, 22039, 19606, 14336, 10976, 
    8616, 3033, -2636, -5473, -9695, -14545, -17433, -20609, -23240, -26171, 
    -28552, -29454, -29689, -30081, -30902, -28600, -27230, -24815, -21503, 
    -19895, -15244, -11718, -6762, -3960, 1596, 4960, 8252, 13102, 17429, 
    20268, 22995, 24844, 27302, 30590, 30736, 31109, 30788, 29267, 26566, 
    24378, 22851, 20449, 16055, 11683, 6662, 2409, -820, -3768, -8614, 
    -13640, -18009, -20940, -22948, -26667, -28205, -30405, -30146, -30645, 
    -30111, -29407, -26135, -24723, -22028, -19284, -16944, -13346, -8658, 
    -4325, 991, 5800, 10089, 13638, 16223, 19167, 23302, 25287, 28218, 29044, 
    29967, 30671, 30070, 30203, 28006, 26056, 23199, 20414, 15705, 12740, 
    7358, 3684, -561, -5277, -9428, -11812, -17448, -21059, -23518, -26612, 
    -29267, -29241, -29616, -30438, -28946, -28970, -28568, -25505, -22516, 
    -20820, -15443, -12554, -8245, -5246, -212, 4145, 7795, 13614, 16723, 
    19936, 21693, 26239, 28188, 28893, 29745, 31170, 30613, 30141, 27717, 
    26247, 21780, 19421, 16672, 12121, 8811, 4500, -466, -5698, -8572, 
    -11913, -15907, -19973, -23025, -25149, -26702, -29673, -30528, -31870, 
    -29362, -28801, -27993, -25706, -24180, -20363, -16438, -13918, -9452, 
    -4623, -1755, 3325, 9267, 11721, 16598, 19058, 23745, 25960, 27817, 
    28853, 29401, 30020, 30336, 29852, 28943, 27433, 24228, 20601, 17321, 
    12110, 10002, 5341, 191, -3836, -8195, -10937, -16180, -19945, -24549, 
    -26636, -28321, -29557, -30375, -30788, -31597, -29575, -28752, -27405, 
    -24113, -22293, -17797, -12797, -10145, -5123, -676, 2860, 6574, 10957, 
    16439, 19037, 22116, 23975, 26508, 29378, 31363, 30144, 29096, 29026, 
    28283, 25811, 23273, 22733, 18588, 13912, 10824, 6325, -161, -2642, 
    -7838, -10513, -15113, -19245, -21518, -25369, -28220, -28736, -29888, 
    -29884, -30459, -28744, -28483, -25824, -24670, -21097, -18718, -13627, 
    -11057, -5003, -1908, 2063, 6408, 12775, 15488, 18865, 21632, 25403, 
    26414, 29467, 29812, 31182, 31188, 31364, 28175, 28235, 25068, 21892, 
    17512, 13708, 9762, 5458, 2210, -2930, -6283, -10375, -14938, -19012, 
    -22423, -25806, -27371, -29566, -30059, -31208, -31523, -30283, -30190, 
    -26611, -25880, -20371, -17716, -13668, -11561, -6904, -2189, 3140, 7561, 
    10712, 14609, 19574, 23105, 25369, 26200, 28801, 29944, 29923, 29866, 
    31633, 29421, 27902, 24467, 20400, 19686, 15736, 10751, 6130, 2105, 
    -1482, -5867, -12066, -13732, -18916, -21581, -24387, -27454, -30152, 
    -31564, -31123, -30891, -29695, -27598, -28635, -26083, -23128, -18852, 
    -16421, -9858, -7676, -1629, 2172, 7076, 10743, 14918, 17625, 22169, 
    25963, 25974, 29406, 31787, 29985, 30278, 31419, 29090, 28086, 24544, 
    21670, 18211, 13785, 10140, 6613, 1719, -1295, -7536, -9510, -13843, 
    -19146, -20926, -22939, -27150, -29747, -28866, -29321, -30423, -28621, 
    -29852, -26721, -25017, -22633, -19033, -16365, -11388, -8167, -2197, 
    963, 5912, 10353, 15913, 17258, 21279, 23556, 25925, 29038, 30980, 29621, 
    31054, 31067, 29579, 26571, 24525, 20686, 18780, 14952, 10368, 6570, 
    3208, -2877, -4460, -9213, -15250, -19005, -21187, -25076, -26673, 
    -26856, -30057, -30591, -30127, -30514, -30346, -28436, -25451, -22843, 
    -19107, -15283, -12481, -7903, -2763, 2864, 6347, 10148, 13114, 17077, 
    21765, 22849, 26368, 29650, 30777, 30417, 30705, 28904, 27748, 26758, 
    24714, 21220, 19609, 16278, 11794, 7272, 2679, -1879, -5274, -10148, 
    -13301, -17921, -21327, -23380, -25024, -27527, -30547, -29531, -30757, 
    -30966, -28511, -26700, -25564, -22424, -19906, -15748, -11713, -6115, 
    -4383, 348, 5007, 9438, 14668, 17541, 21236, 23227, 25414, 27863, 30203, 
    29957, 31593, 31638, 28863, 28889, 25123, 23377, 19994, 15875, 11781, 
    7398, 3145, -782, -5336, -9392, -12494, -16957, -22354, -23969, -25505, 
    -26949, -28049, -28850, -31069, -29909, -28772, -27274, -25437, -22564, 
    -20701, -17032, -11989, -7126, -2449, 945, 4850, 9104, 12754, 18246, 
    20208, 24049, 27788, 28287, 29239, 29561, 29804, 29289, 30860, 28534, 
    25531, 22346, 18704, 17737, 13050, 8113, 3671, 273, -5119, -8234, -11572, 
    -16904, -19952, -24928, -26168, -26495, -30274, -30876, -29439, -30674, 
    -28322, -28164, -26247, -23631, -20112, -15400, -11507, -8733, -4574, 
    240, 3329, 8156, 12806, 16663, 20491, 23636, 25936, 27198, 29626, 29852, 
    29786, 29894, 29536, 28218, 27043, 24146, 19637, 16638, 14022, 9849, 
    5516, 540, -5758, -7138, -12433, -16873, -20939, -24373, -24350, -27939, 
    -30084, -29606, -29863, -29847, -28697, -28640, -26064, -24229, -19421, 
    -16551, -14596, -8576, -4304, -927, 3416, 7566, 13684, 16113, 19183, 
    21653, 25404, 28770, 29348, 31695, 29376, 31506, 29068, 29104, 27281, 
    23954, 21447, 17519, 12308, 10569, 6150, -905, -3142, -6982, -12048, 
    -15320, -19364, -23167, -25596, -28159, -29695, -30423, -30950, -30913, 
    -30373, -29055, -27781, -24657, -20561, -17426, -11966, -10981, -5800, 
    -1126, 2726, 7807, 12588, 15752, 19680, 22958, 24952, 27779, 30250, 
    30800, 31534, 30670, 30662, 28032, 26793, 24764, 22242, 17464, 13528, 
    9356, 4416, 2570, -3871, -6931, -12346, -15424, -19768, -22289, -25832, 
    -27921, -28469, -29491, -29005, -31183, -29767, -29186, -28124, -25006, 
    -20688, -17692, -13923, -9028, -6279, -1535, 3569, 7822, 11462, 15638, 
    18879, 23453, 25407, 28750, 29601, 29337, 30329, 30382, 30460, 29636, 
    25230, 24480, 19898, 18293, 14377, 9531, 5226, 1297, -2846, -8608, 
    -11128, -15421, -18148, -22646, -25158, -27562, -30610, -30565, -31312, 
    -30584, -28390, -28999, -28489, -23755, -20861, -18072, -14081, -9868, 
    -6145, -1855, 3060, 7416, 11247, 15465, 19157, 20736, 26324, 27689, 
    28671, 29578, 29472, 30083, 30534, 28788, 26780, 25812, 21613, 19213, 
    14359, 11569, 6280, 1337, -2118, -5206, -11009, -14967, -18418, -23413, 
    -24593, -27027, -30012, -31190, -29088, -31223, -28886, -29924, -26860, 
    -24602, -23525, -19185, -13833, -11921, -5992, -2545, 2179, 7205, 9507, 
    14760, 18479, 22316, 26059, 26374, 29177, 30934, 31225, 30724, 29977, 
    27568, 27599, 24341, 21874, 18736, 15392, 9393, 5675, 1583, -1111, -6074, 
    -11304, -14208, -18216, -20856, -23344, -26408, -28666, -30758, -31190, 
    -29656, -31560, -28815, -25757, -26325, -22724, -18912, -14260, -9789, 
    -6046, -1716, 758, 6144, 11211, 12599, 17536, 22240, 25254, 26729, 29213, 
    30397, 30646, 31553, 29111, 28414, 28043, 25223, 20751, 18022, 15067, 
    11480, 7071, 1513, -911, -5423, -10156, -13342, -16630, -21269, -24305, 
    -26952, -28312, -29345, -30255, -31021, -29433, -27959, -27032, -24759, 
    -22007, -19977, -14343, -11305, -8025, -2205, 1668, 6341, 9858, 14600, 
    16640, 21943, 23993, 26629, 28441, 30267, 30719, 30320, 31263, 28731, 
    28850, 26392, 22277, 17921, 14983, 12866, 8844, 4522, -1279, -3986, 
    -10994, -14606, -16531, -19384, -22569, -26743, -28419, -28972, -31539, 
    -30622, -31011, -28078, -27211, -26934, -23652, -20523, -15512, -12317, 
    -7791, -3620, 952, 5725, 10862, 14178, 18011, 21464, 24314, 24976, 26938, 
    29841, 31743, 30752, 30446, 30567, 26846, 26533, 22616, 19410, 15011, 
    11386, 8291, 3312, -2032, -3973, -8154, -13098, -17706, -20049, -23574, 
    -26569, -28550, -31457, -31715, -29046, -29108, -29593, -26868, -24888, 
    -22280, -18755, -15015, -12758, -9834, -4567, 769, 5768, 9781, 12172, 
    15870, 21814, 24441, 26257, 27474, 30243, 29962, 32079, 31606, 30362, 
    27655, 24777, 23019, 19669, 16748, 11754, 9235, 3648, -1024, -4490, 
    -7913, -11387, -16292, -21500, -24799, -26579, -29237, -30933, -29223, 
    -30248, -30415, -30478, -26919, -26319, -24217, -21997, -17243, -13785, 
    -7281, -3414, 481, 3183, 8903, 12670, 17177, 21055, 22276, 27141, 29499, 
    30952, 31233, 29695, 31504, 29583, 28767, 25777, 22845, 21261, 16803, 
    13611, 9711, 4890, -389, -5241, -9238, -13250, -16360, -18578, -23228, 
    -25339, -27557, -30178, -31258, -30436, -29178, -28486, -27316, -25477, 
    -24572, -19275, -16427, -13449, -9029, -5400, -1085, 4464, 8085, 12526, 
    17176, 19600, 24208, 23965, 28503, 27839, 29233, 30921, 30205, 29351, 
    29332, 26772, 23781, 21396, 17075, 12701, 8603, 5274, 2296, -4857, -8318, 
    -12048, -14780, -18061, -21347, -25245, -28703, -30198, -30124, -30742, 
    -29964, -29712, -28206, -27018, -23694, -20470, -16707, -12566, -9067, 
    -4932, -1916, 4921, 6791, 11743, 15241, 19187, 24308, 25566, 28474, 
    30111, 31793, 29441, 30431, 30380, 29749, 25570, 23831, 22094, 17054, 
    15152, 9845, 4801, 949, -3629, -9425, -12654, -15723, -19543, -21954, 
    -24765, -26953, -30046, -30602, -30952, -30094, -30411, -27655, -27591, 
    -24655, -22119, -17734, -15261, -10673, -5315, -1352, 4218, 7548, 11747, 
    14732, 19437, 21884, 26748, 26676, 30147, 30341, 31745, 30589, 28566, 
    28832, 26076, 24452, 20415, 19245, 14359, 10605, 5658, 498, -2815, -7093, 
    -11072, -14545, -18121, -23487, -24834, -26014, -29043, -31179, -31495, 
    -29766, -30396, -27646, -27052, -25407, -22278, -18238, -14422, -10332, 
    -5918, -3166, 3872, 7289, 11201, 16495, 17815, 23027, 24035, 27073, 
    29197, 29148, 30590, 30920, 29520, 28251, 25876, 25511, 21539, 18542, 
    14008, 10332, 6357, 2874, -2505, -7680, -11496, -15204, -17349, -21632, 
    -24016, -26797, -27559, -31012, -32034, -29069, -29460, -28907, -26568, 
    -25019, -22260, -18132, -14591, -11241, -7322, -1647, 2356, 5686, 11053, 
    13844, 16860, 22219, 25098, 28030, 29571, 31298, 30482, 29448, 31506, 
    28730, 26615, 25618, 22200, 18357, 15646, 11576, 7026, 2222, -1904, 
    -6684, -10809, -15129, -19293, -21155, -23905, -25394, -30210, -29609, 
    -30537, -31303, -30075, -28157, -27214, -26522, -23046, -17226, -14518, 
    -10123, -7244, -1201, 1377, 5222, 11351, 14261, 19293, 20374, 24656, 
    26999, 30221, 30033, 31822, 31041, 29297, 27675, 28384, 23891, 20835, 
    19017, 15481, 12525, 6451, 2960, -2057, -5438, -8831, -13882, -17070, 
    -21016, -25279, -27085, -28179, -28936, -30612, -31250, -30884, -29458, 
    -27079, -24674, -22172, -18308, -15464, -11735, -6640, -3389, 1934, 4955, 
    9485, 13953, 16781, 22992, 22652, 26667, 27658, 28739, 32084, 30723, 
    31121, 29968, 27475, 27089, 23380, 19314, 16232, 10726, 8349, 2357, 
    -1267, -4962, -9337, -14541, -18924, -21325, -22806, -25875, -28644, 
    -30193, -31832, -31117, -30399, -28814, -26688, -25334, -22755, -19054, 
    -16384, -12746, -6608, -4192, 1842, 5458, 9618, 12758, 17120, 20305, 
    22512, 25070, 28060, 29364, 30381, 31493, 30450, 29071, 27276, 25143, 
    21358, 19478, 17129, 12151, 7714, 3729, -747, -6118, -9898, -13909, 
    -18409, -19146, -23549, -27229, -28357, -29117, -30272, -31732, -31160, 
    -30400, -27080, -24482, -23585, -18020, -15444, -13325, -7695, -3410, 
    559, 5475, 10249, 14947, 16480, 21352, 23073, 24664, 27792, 30072, 31554, 
    30541, 31686, 30430, 27282, 24513, 23891, 19814, 15079, 12573, 7774, 
    3886, 944, -6395, -9694, -12645, -15555, -20323, -23205, -26646, -28498, 
    -29259, -31180, -30031, -30809, -30187, -28411, -26613, -23301, -21130, 
    -15874, -13671, -9701, -4809, -389, 3961, 8786, 12040, 17821, 19580, 
    23643, 25346, 28422, 30161, 30335, 30271, 30701, 29688, 27196, 24710, 
    23174, 20761, 17011, 13412, 9270, 3406, -665, -4915, -8122, -12259, 
    -15221, -18748, -23638, -25593, -26708, -30506, -31052, -30638, -31114, 
    -29231, -29014, -26686, -23102, -19490, -16811, -12963, -10029, -3200, 
    -1335, 5495, 7575, 11813, 15806, 20109, 22751, 24785, 27921, 28698, 
    29999, 29372, 29840, 29285, 28571, 25404, 23567, 20553, 18701, 13818, 
    8935, 4774, 289, -4070, -9671, -12621, -16204, -18886, -23704, -24638, 
    -27099, -27779, -29338, -30737, -29998, -28018, -28854, -25579, -24129, 
    -20170, -18172, -14614, -10286, -4986, -1115, 3827, 7776, 12359, 14219, 
    19900, 22210, 26022, 26950, 28475, 31401, 30919, 31077, 31238, 28205, 
    25292, 23576, 20145, 18074, 13896, 11121, 6137, 750, -3859, -6018, 
    -11885, -14449, -19906, -24141, -26770, -27415, -27723, -30908, -30676, 
    -31550, -29060, -27634, -26637, -23374, -21093, -18298, -14562, -11708, 
    -6479, -28, 3838, 8595, 10681, 15737, 18513, 21019, 25150, 28804, 27823, 
    29274, 30548, 30630, 29441, 28554, 28246, 24567, 21827, 18335, 13564, 
    11721, 6235, 127, -2530, -7154, -10770, -14507, -19732, -23253, -23729, 
    -26127, -28954, -31534, -31468, -29303, -30247, -29203, -26833, -25636, 
    -21429, -17869, -15254, -9146, -5722, -1336, 2158, 6022, 12721, 15068, 
    18674, 22351, 23794, 27217, 29435, 31380, 31350, 30564, 30646, 30139, 
    27599, 23407, 21544, 18916, 14813, 10742, 6915, 1456, -3567, -4989, 
    -11534, -14275, -19588, -20836, -25555, -26126, -28055, -31047, -30826, 
    -30822, -30371, -28977, -27872, -24848, -22702, -18495, -14907, -10772, 
    -7035, -1599, 2325, 6622, 9868, 14951, 18570, 22578, 25533, 28673, 29271, 
    30527, 31062, 30502, 30236, 27385, 26868, 24103, 22071, 19572, 13778, 
    10823, 5428, 2371, -1747, -5475, -9621, -15495, -17357, -20656, -24566, 
    -27237, -29946, -29495, -31343, -30290, -29291, -29043, -26398, -24789, 
    -22668, -19857, -16646, -11662, -6599, -2871, 2213, 5889, 11357, 14445, 
    17282, 23130, 24072, 27583, 30233, 28578, 32117, 30476, 30276, 27268, 
    26962, 25594, 22406, 18148, 15624, 11337, 7623, 3078, -2750, -6776, 
    -11085, -13342, -16984, -21747, -23946, -26980, -27651, -29620, -31684, 
    -30178, -30526, -28487, -26061, -25272, -23245, -19251, -16776, -10585, 
    -7688, -2037, 433, 4943, 10081, 14225, 17758, 20485, 23972, 27609, 28155, 
    30805, 29806, 29443, 29881, 30579, 28430, 26571, 22228, 19520, 15915, 
    11765, 7617, 2165, -501, -5151, -9675, -13728, -18926, -21858, -24063, 
    -27688, -29175, -30101, -31830, -32305, -28788, -29757, -26762, -26315, 
    -23393, -19416, -16847, -11770, -9178, -3997, 292, 5398, 10115, 13623, 
    17677, 20959, 23962, 25589, 28392, 30069, 31062, 31055, 28685, 28220, 
    27422, 23977, 23903, 20729, 16486, 10665, 7792, 3624, 330, -5198, -9115, 
    -12210, -16913, -21390, -22884, -26560, -28532, -30948, -29146, -31321, 
    -31052, -28019, -26024, -25041, -22189, -19349, -16785, -13514, -8138, 
    -4218, 1607, 3717, 11017, 13017, 17280, 19978, 23085, 26075, 28900, 
    31302, 30004, 31476, 29830, 30077, 28630, 26553, 22360, 18958, 17498, 
    11955, 9160, 3904, -1755, -3392, -8925, -14194, -16582, -20031, -22699, 
    -25691, -27764, -29650, -30425, -30062, -29498, -30156, -26699, -26648, 
    -22411, -21149, -16259, -12858, -8746, -4795, -178, 4532, 9098, 11831, 
    15088, 19804, 24422, 26207, 28074, 28864, 31573, 30021, 30825, 29255, 
    28608, 25170, 23641, 20950, 16789, 13194, 8990, 5736, 568, -5117, -8251, 
    -10935, -17669, -19728, -23719, -25062, -26436, -29493, -29477, -30110, 
    -31328, -29533, -29590, -26722, -22916, -19863, -16572, -12673, -8365, 
    -5778, 149, 4334, 7961, 13847, 16719, 19503, 22777, 25408, 28236, 30073, 
    29988, 31539, 29432, 29982, 27745, 26788, 22125, 20870, 16500, 12833, 
    9654, 6172, 1452, -3344, -6248, -12376, -16111, -20348, -24019, -25750, 
    -27126, -28906, -29885, -30641, -28811, -29873, -28534, -27066, -25133, 
    -21016, -19096, -13680, -9369, -4711, 182, 3791, 7152, 12570, 16009, 
    18070, 21029, 26778, 26964, 27707, 31416, 30821, 29104, 30301, 28162, 
    25738, 23933, 20412, 17581, 15026, 9455, 5528, 124, -2488, -8844, -10518, 
    -14426, -17791, -21877, -23884, -27835, -28800, -31322, -29667, -30048, 
    -30711, -27317, -26777, -24478, -21719, -18419, -14757, -10085, -6401, 
    -819, 4083, 7825, 11115, 14531, 18993, 22674, 26364, 27361, 28370, 31453, 
    31506, 30306, 29566, 29173, 25063, 25146, 21224, 17660, 14525, 10486, 6124, 
    1239, -3871, -6758, -11274, -15074, -18117, -22506, -26510, -26515, 
    -28731, -29967, -31624, -31938, -30839, -27950, -27366, -25586, -21394, 
    -17325, -13693, -11753, -5961, -2807, 2714, 6254, 12439, 15348, 18796, 
    21951, 25268, 28424, 29859, 30990, 31458, 31075, 29606, 28073, 26267, 
    24500, 20737, 18178, 14116, 12378, 6655, 1100, -3340, -6551, -10482, 
    -14305, -17194, -21944, -25125, -28053, -29361, -29114, -32114, -30553, 
    -30305, -29126, -26752, -24988, -21333, -18936, -14294, -10442, -5375, 
    -2457, 2458, 6308, 11032, 14352, 18403, 22609, 25708, 26572, 29146, 
    30221, 30975, 30996, 29581, 30200, 26350, 23962, 21106, 17416, 14385, 
    9477, 5791, 2546, -1030, -5759, -11186, -13992, -19684, -20574, -26114, 
    -26448, -29604, -30835, -30329, -30036, -30939, -29057, -27319, -25366, 
    -20864, -19360, -14516, -10810, -7220, -2797, 2328, 6150, 9400, 14423, 
    18487, 21229, 24657, 28361, 29849, 29928, 30811, 30772, 30061, 29309, 
    26031, 24904, 22116, 18582, 16576, 12768, 7221, 4109, -1890, -5451, 
    -10330, -14502, -19657, -21609, -23329, -26354, -28118, -30077, -30327, 
    -30638, -29599, -28812, -26960, -25032, -21766, -20239, -16474, -11224, 
    -6949, -1960, 1652, 5864, 10719, 13837, 16253, 21151, 24484, 25773, 
    27864, 28400, 31632, 31346, 30799, 28315, 27752, 25764, 23327, 17997, 
    15259, 11093, 8687, 2266, -1168, -3828, -9236, -13899, -16667, -20307, 
    -23652, -26256, -29186, -30618, -31094, -30816, -31325, -28340, -28129, 
    -25381, -21514, -18474, -15558, -12664, -8961, -3798, -205, 4846, 11032, 
    13651, 17313, 20641, 23686, 25445, 27583, 29523, 29119, 30567, 29958, 
    28429, 27371, 25033, 21844, 19976, 17729, 11547, 8011, 2933, -1442, 
    -3942, -9050, -13458, -16782, -20912, -22498, -25427, -29643, -30420, 
    -30752, -29835, -29969, -28835, -27919, -25230, -22549, -19746, -15294, 
    -12570, -8185, -3719, -740, 6493, 8416, 12904, 17888, 21950, 22664, 
    26889, 26559, 30967, 31900, 31039, 30616, 29478, 28697, 25689, 23194, 
    20145, 16248, 11381, 6690, 3325, 919, -6310, -8590, -11991, -16578, 
    -21032, -22566, -25558, -29607, -28828, -31192, -30850, -30084, -29741, 
    -28069, -25357, -24558, -21448, -17427, -12790, -7138, -4152, -1386, 
    4927, 7809, 11119, 17653, 20470, 23192, 25471, 26870, 29337, 30406, 
    30001, 31260, 29735, 28387, 25583, 24529, 19369, 16201, 14100, 9118, 
    4419, -306, -3993, -8527, -12336, -16804, -19812, -21987, -25092, -28159, 
    -28457, -31568, -30871, -30467, -30121, -27955, -27701, -23057, -19401, 
    -16387, -12459, -10128, -5249, 437, 4262, 7843, 12282, 16529, 18647, 
    23520, 26587, 28510, 28775, 29378, 30087, 29368, 29161, 29494, 26723, 
    22591, 19697, 17083, 14000, 9673, 3505, 1108, -3407, -8269, -10837, 
    -17069, -18841, -22381, -23767, -29214, -29749, -30055, -32586, -29534, 
    -30547, -27811, -25308, -24018, -20899, -17543, -13017, -10195, -5764, 
    -606, 4330, 8570, 10815, 16812, 19989, 22695, 26299, 28140, 29612, 31308, 
    30164, 32308, 30197, 29278, 26617, 25084, 21757, 18295, 13252, 10403, 
    5672, 943, -2866, -7222, -12573, -14928, -19639, -23805, -25691, -26498, 
    -28002, -31893, -31413, -29269, -31557, -28519, -25850, -23984, -21312, 
    -17099, -14015, -11493, -6402, -1064, 3460, 7043, 12060, 15134, 18692, 
    22455, 24531, 27053, 30135, 31041, 31254, 30810, 30323, 27918, 26598, 
    24639, 21686, 18612, 15168, 11018, 5664, 1988, -2724, -6539, -10139, 
    -15156, -17754, -22122, -25430, -25959, -28345, -28796, -30245, -31849, 
    -30649, -29956, -25038, -23733, -21990, -17436, -15211, -9425, -5835, 
    -1612, 2651, 6021, 11469, 15270, 17943, 22828, 26117, 26994, 27887, 
    29339, 30275, 30251, 29662, 28927, 28026, 24758, 21157, 19040, 15045, 
    10058, 6182, 1855, -2361, -5515, -11515, -14239, -18722, -22410, -25658, 
    -27824, -30120, -31306, -29408, -30965, -29523, -29828, -27219, -24907, 
    -21433, -19622, -13350, -10121, -6954, -1020, 1539, 6631, 10222, 15232, 
    18569, 21091, 23873, 27452, 30191, 28459, 30827, 30948, 30312, 27477, 
    27980, 24469, 21392, 19394, 13849, 11414, 6539, 1667, -1587, -6256, 
    -12055, -14518, -17578, -21760, -24207, -26647, -29223, -29723, -30719, 
    -30798, -30089, -28814, -27552, -25212, -20568, -18370, -14959, -11528, 
    -8043, -2287, 1629, 6377, 8984, 15234, 16934, 19999, 23931, 26337, 29193, 
    29200, 32075, 29308, 29397, 29273, 26146, 25804, 22490, 18226, 13927, 
    12853, 8319, 2616, -2491, -5220, -9707, -13541, -19685, -21707, -24926, 
    -25445, -28737, -31315, -30368, -30531, -29063, -28432, -25780, -25744, 
    -22671, -18827, -16584, -12210, -8049, -3685, 1257, 6389, 10907, 13514, 
    17881, 21912, 23957, 27951, 28916, 29386, 30776, 32129, 29096, 30124, 
    27311, 25251, 22311, 20084, 16145, 13516, 8901, 3983, -149, -6617, -9073, 
    -13343, -17313, -21727, -23752, -25057, -28637, -30009, -29763, -30697, 
    -28577, -29368, -26894, -25204, -22116, -18911, -16632, -12852, -8453, 
    -3902, -188, 4572, 8576, 13342, 16116, 20479, 23920, 27155, 27105, 29662, 
    30581, 29584, 30637, 29972, 27844, 26111, 22612, 18940, 16589, 13131, 
    8092, 2590, 944, -5214, -8459, -12713, -17288, -20966, -24436, -27586, 
    -27667, -29027, -31343, -32268, -31733, -28384, -28657, -24324, -22760, 
    -19289, -16017, -12403, -7839, -3811, -499, 3821, 9354, 13980, 15950, 
    21002, 24700, 26088, 27700, 29078, 29493, 31860, 29770, 28969, 26939, 
    25073, 23051, 20014, 16336, 10770, 8446, 3454, 1034, -4602, -8777, 
    -13563, -16597, -20490, -23629, -26730, -27625, -29006, -30949, -32312, 
    -30857, -29288, -29063, -26872, -23775, -20281, -17352, -12516, -8634, 
    -4786, -1128, 4194, 9710, 12820, 17527, 21447, 22342, 25119, 29491, 
    29886, 30128, 31457, 31168, 28881, 27675, 27487, 24422, 20289, 15224, 
    12799, 9257, 4676, -649, -2900, -7414, -12217, -15447, -20159, -23707, 
    -25805, -26501, -28326, -30151, -29885, -31236, -31056, -28442, -25622, 
    -23466, -21176, -16869, -14665, -8760, -3669, -557, 4343, 7924, 12880, 
    16187, 20169, 21243, 25006, 27894, 30227, 32027, 31080, 31262, 30137, 
    27847, 25206, 23633, 21584, 18735, 13168, 9814, 5177, -456, -2277, -8097, 
    -12588, -15233, -19896, -22709, -25161, -27622, -29677, -31560, -30438, 
    -30640, -30100, -28181, -27649, -23567, -21974, -18169, -11928, -9342, 
    -5676, -1750, 2415, 6593, 12298, 16851, 19261, 21604, 26600, 27907, 
    29901, 31242, 30225, 31664, 30317, 27816, 26421, 25676, 19824, 19113, 
    14015, 8236, 4153, 989, -3418, -7960, -12613, -15069, -19483, -24244, 
    -25614, -27915, -29679, -30722, -31290, -30415, -28793, -29908, -25724, 
    -24297, -21728, -19293, -14318, -11223, -4771, -656, 2346, 6878, 10858, 
    16869, 19662, 21927, 24234, 27414, 27901, 29168, 30737, 30759, 29941, 
    28173, 26703, 24040, 21017, 16823, 14689, 11536, 5899, 1311, -2405, 
    -6439, -12554, -14635, -18852, -22577, -24627, -28037, -30344, -29900, 
    -30902, -29581, -30896, -29348, -26523, -23812, -21274, -17736, -14297, 
    -10032, -7282, -2410, 2136, 6150, 10183, 15559, 17705, 21041, 23908, 
    27231, 29158, 29198, 30193, 30321, 29996, 28822, 26217, 25307, 21793, 
    18190, 13876, 10161, 6641, 343, -1695, -6906, -12133, -15534, -18864, 
    -21273, -24597, -27442, -29641, -29003, -30874, -31067, -29714, -30094, 
    -26886, -23946, -22532, -17896, -15039, -11180, -5453, -3044, 3048, 6808, 
    9557, 15500, 18668, 21575, 24046, 27046, 29450, 29043, 30358, 30024, 
    30910, 27611, 26990, 24706, 20512, 17027, 15162, 10405, 8095, 3600, 
    -2149, -7122, -10093, -15413, -18673, -23152, -24163, -27709, -28100, 
    -28675, -30637, -30950, -31702, -28711, -27442, -24798, -22490, -19600, 
    -16363, -10327, -5924, -2766, 816, 7126, 10983, 13628, 18766, 21288, 24925, 
    26716, 28946, 30033, 31563, 29194, 31063, 28175, 27778, 23913, 22092, 
    20446, 14588, 9924, 7220, 1951, -1376, -5713, -10076, -14182, -17481, 
    -20744, -23600, -26621, -28142, -29970, -30422, -29558, -30017, -29480, 
    -27333, -25631, -21262, -18737, -16725, -11305, -8151, -2238, 1616, 5221, 
    10152, 13198, 17725, 21406, 24016, 27061, 27798, 30388, 30461, 30060, 
    30617, 27872, 28138, 25055, 22897, 19793, 16874, 11679, 6856, 3273, -343, 
    -5255, -9482, -12982, -16762, -22206, -22906, -28312, -28029, -30635, 
    -30809, -29434, -31068, -28526, -27159, -26246, -22865, -18126, -15697, 
    -13402, -8584, -3242, 671, 6408, 10238, 13915, 17288, 20872, 22493, 
    26307, 27059, 29672, 30917, 30778, 29042, 30487, 28147, 26180, 22349, 
    19380, 16200, 12091, 8397, 3383, -737, -4176, -8271, -13617, -17159, 
    -19417, -24298, -26653, -29951, -29651, -30842, -31881, -30970, -29545, 
    -26604, -26909, -22863, -19414, -14989, -12733, -7269, -3971, -813, 4819, 
    8013, 13223, 17277, 19813, 23492, 25744, 27188, 28863, 29148, 31582, 
    29936, 29299, 27620, 25930, 24343, 20055, 17275, 14016, 9802, 5050, -898, 
    -4718, -8522, -12645, -15848, -20705, -23487, -26088, -27174, -30305, 
    -30492, -30071, -29464, -30846, -28363, -24874, -23741, -21311, -16047, 
    -13844, -9109, -4550, -543, 3395, 8613, 12924, 17005, 20594, 22106, 
    25180, 27995, 29951, 29470, 30731, 29797, 30487, 26808, 25824, 24573, 
    21694, 17085, 11968, 8940, 5451, 16, -3841, -6704, -11507, -16061, 
    -19917, -22870, -25990, -26693, -30177, -29740, -29865, -30665, -28424, 
    -27010, -25004, -23508, -20232, -16239, -12621, -10061, -3319, -528, 
    4255, 8737, 11752, 16208, 18667, 22095, 25711, 28116, 29201, 32333, 
    31630, 31586, 31341, 28524, 26191, 24568, 21341, 17233, 13851, 10367, 
    4500, 1272, -4100, -7801, -13538, -15715, -18444, -23778, -24974, -27656, 
    -30998, -30078, -30299, -30740, -29257, -27518, -25584, -24260, -21161, 
    -17127, -14670, -9088, -5250, -1298, 4375, 8496, 11005, 15478, 20127, 
    22970, 26123, 27886, 29385, 31620, 31964, 30590, 31015, 28139, 27464, 
    23878, 20571, 18304, 13561, 8248, 4926, 1206, -3603, -6911, -11745, 
    -15964, -20537, -21191, -23725, -27468, -29598, -30658, -31772, -31299, 
    -30101, -29257, -26047, -25664, -19834, -17744, -13392, -10879, -5604, 
    -2426, 2502, 7250, 11970, 14279, 19928, 22132, 26632, 27830, 30141, 
    28932, 29868, 30901, 29161, 28366, 25150, 25374, 20700, 17645, 15602, 
    9662, 4086, 3283, -3955, -6292, -10105, -14676, -19379, -22238, -24446, 
    -26474, -28768, -30781, -29165, -29977, -31724, -29937, -25415, -22810, 
    -22351, -18017, -15162, -9610, -5154, -1614, 3569, 6710, 12839, 16243, 
    18488, 22363, 26285, 26668, 27553, 31832, 31513, 32234, 29883, 28270, 
    27652, 24508, 21417, 18281, 14522, 10721, 6676, 2189, -3136, -7621, 
    -12317, -14014, -18635, -22445, -24941, -27255, -29154, -28964, -30716, 
    -30919, -30350, -28079, -27098, -24001, -20549, -18822, -14472, -10133, 
    -6468, -2017, 3242, 7738, 10957, 14550, 18349, 21327, 25706, 26624, 
    28813, 30246, 29089, 29912, 29665, 29310, 26933, 23366, 22794, 17968, 
    14655, 11127, 5860, 2497, -2460, -6715, -9090, -14901, -19491, -21312, 
    -24868, -26676, -27489, -30276, -30733, -30494, -28990, -27916, -26667, 
    -24311, -22305, -18630, -16217, -10765, -6785, -2580, 1111, 6661, 10445, 
    15694, 16491, 21970, 23523, 26586, 29453, 30664, 30757, 31796, 30091, 
    29196, 27038, 24781, 20987, 19091, 14413, 10701, 6664, 3802, -445, -4251, 
    -8688, -15835, -17920, -20922, -24680, -27817, -28907, -28883, -29447, 
    -30706, -29839, -29241, -27321, -26285, -22063, -18400, -15685, -11846, 
    -6933, -4391, 1734, 4688, 9876, 14157, 17514, 21060, 23981, 26409, 28981, 
    29616, 29866, 30077, 30615, 28918, 27379, 24036, 22895, 18662, 17292, 
    11300, 6131, 4808, -735, -5332, -9628, -14165, -17956, -21112, -25068, 
    -27159, -28642, -29973, -30002, -31699, -31037, -29391, -26700, -26135, 
    -22375, -21157, -15983, -13106, -7116, -1984, 1595, 5212, 8916, 13277, 
    17210, 20568, 24632, 26890, 28511, 29421, 30057, 30858, 30598, 29522, 
    26965, 25341, 23398, 19201, 15186, 12386, 7978, 3032, -1107, -3985, 
    -8882, -13661, -18259, -20979, -23001, -25548, -29205, -31330, -30142, 
    -32545, -29757, -29615, -27491, -25685, -22896, -20362, -14833, -11523, 
    -9033, -4286, -1095, 4759, 8641, 14504, 16714, 19100, 22956, 25342, 
    27940, 30126, 29072, 30799, 30826, 28428, 28105, 24766, 22920, 19713, 
    15912, 13910, 9551, 3746, -428, -3119, -8584, -13140, -16662, -18932, 
    -23789, -26067, -28885, -30660, -29896, -30546, -31603, -28313, -29105, 
    -25380, -23463, -19881, -17134, -13277, -8748, -3545, -988, 4848, 9425, 
    11997, 16760, 20372, 22528, 24293, 28440, 30656, 31203, 30180, 30682, 
    30797, 28000, 25762, 23138, 19764, 15837, 12842, 9668, 3183, -294, -3898, 
    -7712, -11129, -17124, -20991, -22548, -26537, -28241, -29546, -30045, 
    -30768, -31333, -30308, -29523, -27490, -23783, -19461, -16915, -13143, 
    -9495, -5044, -97, 3943, 8343, 12038, 17271, 19791, 23118, 26101, 26710, 
    29529, 30121, 29939, 30649, 29334, 27302, 26961, 22194, 21138, 16717, 
    12867, 8222, 6217, 657, -3336, -7833, -12956, -17773, -18486, -23084, 
    -24195, -27346, -30062, -31075, -30773, -31024, -29411, -27670, -26180, 
    -23595, -22053, -16679, -13244, -9698, -6708, -1400, 2484, 7758, 11104, 
    14504, 19725, 21991, 25128, 28172, 28917, 30104, 30175, 30437, 28278, 
    28499, 26986, 23034, 21235, 18727, 14123, 9160, 6632, 2178, -4079, -7687, 
    -13062, -14938, -18709, -22246, -26650, -27411, -29990, -30678, -31109, 
    -29522, -30331, -28193, -27251, -23317, -22205, -18108, -15080, -10913, 
    -6463, -987, 3599, 7849, 10401, 15242, 19000, 22482, 24706, 28580, 28533, 
    29817, 32048, 30526, 30003, 27974, 26834, 23769, 21519, 18834, 14135, 
    11336, 5797, 1292, -1320, -6019, -10837, -15480, -19696, -22018, -24499, 
    -27074, -30132, -29497, -30746, -31863, -30239, -29228, -25587, -23260, 
    -20201, -19069, -13981, -10701, -6154, -2085, 3558, 6465, 10483, 15467, 
    17481, 20715, 26399, 26245, 28741, 30902, 31404, 31255, 28901, 28956, 
    25956, 25030, 21898, 18406, 14071, 10524, 5564, 2319, -3260, -6857, 
    -11389, -14595, -18536, -22630, -24641, -26929, -28535, -29601, -30765, 
    -29997, -30014, -28166, -25844, -25230, -21122, -18877, -15436, -11549, 
    -6251, -391, 3164, 6231, 11190, 13572, 18204, 20979, 24611, 25991, 27365, 
    30520, 29436, 29519, 30033, 28718, 27538, 25197, 22370, 18673, 14828, 
    12620, 6527, 3113, -1507, -5826, -11268, -14943, -18211, -21997, -23843, 
    -26788, -28791, -29544, -30754, -30647, -30382, -27885, -26716, -24936, 
    -22748, -20172, -14975, -10827, -8812, -2972, 1142, 5636, 9191, 13343, 
    19320, 21467, 25981, 27101, 27643, 28954, 31167, 30482, 30394, 28617, 
    27784, 26781, 22249, 19588, 14545, 11358, 7735, 2174, -2217, -6107, 
    -9917, -15140, -17447, -21481, -25557, -27292, -29404, -29632, -29593, 
    -31189, -30514, -27939, -28979, -26242, -23396, -17657, -15454, -12615, 
    -7316, -2884, 646, 5192, 10556, 12864, 19145, 20919, 23580, 28234, 28232, 
    30905, 31811, 31637, 30751, 28093, 28001, 26784, 22801, 20143, 15365, 
    12202, 7856, 3347, -1371, -5727, -9971, -12366, -18523, -20458, -24166, 
    -26213, -27218, -29915, -30579, -30986, -30982, -29815, -26571, -24815, 
    -22424, -20386, -15695, -12821, -8104, -2938, -249, 5315, 9832, 14301, 
    18796, 20889, 25053, 26048, 28260, 30749, 29831, 31619, 29541, 29847, 
    28737, 26019, 23538, 20148, 16099, 12981, 7808, 4479, -1333, -6720, 
    -8305, -13222, -16158, -21111, -22768, -26851, -29149, -30588, -29603, 
    -29619, -29439, -29089, -27273, -25302, -23211, -20091, -17082, -13907, 
    -9513, -2981, -1073, 5672, 9415, 13796, 16545, 19729, 23898, 26943, 
    28011, 28398, 29826, 30768, 29858, 28992, 27293, 26246, 23892, 19577, 
    18011, 13207, 9011, 5017, -686, -5324, -8958, -12018, -17940, -20093, 
    -24229, -25599, -27423, -30940, -30949, -31422, -30372, -29444, -27253, 
    -25935, -22988, -20270, -17045, -12916, -6787, -5153, 277, 4050, 9319, 
    12202, 17257, 19727, 22752, 25264, 29122, 29136, 29357, 31207, 30431, 
    30845, 28381, 24934, 24365, 21321, 16512, 13161, 9211, 5370, 1816, -4066, 
    -9339, -12334, -16701, -20109, -22729, -25205, -27824, -28804, -30606, 
    -31078, -30089, -29954, -28828, -25038, -22610, -21046, -16654, -13309, 
    -9140, -4113, 433, 4444, 8093, 11791, 16075, 20130, 23134, 25741, 28463, 
    29367, 30561, 30600, 29698, 29407, 29006, 26972, 23341, 19838, 17639, 
    14470, 9488, 5760, 921, -4869, -8276, -12120, -15804, -18663, -23008, 
    -25240, -27867, -30187, -31115, -30784, -29404, -28407, -27665, -26024, 
    -23197, -20058, -16994, -13939, -8684, -4924, 476, 3275, 9089, 12411, 
    14628, 19412, 22490, 26539, 27084, 29074, 29910, 30972, 31351, 30011, 
    30076, 26781, 23104, 20424, 17110, 14352, 9086, 6543, 1310, -2667, -6800, 
    -10662, -14152, -20621, -23140, -24669, -26553, -30251, -29713, -30709, 
    -31243, -29022, -29561, -27389, -23258, -21624, -18016, -14096, -8190, 
    -6466, -172, 2365, 6820, 11098, 15420, 18982, 22402, 25178, 28947, 30195, 
    28846, 31503, 29961, 28758, 28121, 26847, 25670, 21071, 17775, 12972, 
    11473, 6097, 580, -2820, -7463, -12154, -14962, -20151, -21163, -26910, 
    -26861, -27812, -30298, -31581, -30977, -29228, -28885, -26739, -24090, 
    -21113, -17852, -15112, -10430, -6708, -2600, 1950, 7802, 10897, 15701, 
    18666, 22717, 25901, 27524, 28681, 30339, 30538, 31089, 30326, 27848, 
    26626, 24232, 21043, 19362, 14490, 10419, 6000, 2782, -2096, -6355, 
    -10317, -13665, -18148, -22153, -23943, -27037, -28668, -30575, -30006, 
    -30563, -30295, -28289, -27288, -23993, -22845, -18434, -14714, -9968, 
    -6502, -3817, 2939, 8158, 9741, 14469, 19423, 21017, 23217, 26888, 29400, 
    29130, 29070, 30118, 30308, 29004, 26507, 25224, 23144, 17470, 14027, 
    12567, 6014, 2352, -3154, -5061, -10424, -15446, -16801, -22488, -25635, 
    -25986, -28017, -29165, -29798, -29832, -30941, -27834, -27338, -24625, 
    -21555, -19970, -15446, -10701, -6129, -2404, 2882, 5723, 10274, 15096, 
    17871, 21307, 25793, 27339, 29438, 28674, 29851, 31380, 30115, 30200, 
    25454, 25200, 21877, 17596, 15228, 10881, 8272, 2529, -392, -7558, 
    -11016, -14400, -16614, -19847, -23472, -25257, -30337, -29283, -30501, 
    -29945, -29188, -30124, -27723, -26193, -21267, -19761, -14141, -10830, 
    -6179, -2671, 1121, 5823, 9702, 13863, 17749, 20864, 25431, 26068, 28144, 
    28479, 30161, 31852, 29997, 30333, 25949, 24145, 22241, 19564, 14298, 
    10139, 7411, 4132, -1247, -5909, -9402, -13980, -17778, -21763, -24732, 
    -25698, -28855, -29320, -29963, -29547, -30557, -28456, -26151, -25069, 
    -23553, -19301, -15212, -11672, -6996, -3780, -386, 5202, 10569, 13281, 
    17621, 19911, 23872, 27096, 28904, 28422, 29677, 31545, 31313, 29504, 
    28711, 24699, 23038, 20858, 16608, 11075, 7401, 3566, -1336, -5342, 
    -9606, -12952, -18159, -21618, -24957, -26513, -28348, -29440, -31335, 
    -31133, -29527, -30430, -29526, -27441, -22116, -20187, -17217, -13309, 
    -6654, -4904, 1302, 4605, 7712, 13540, 17507, 21067, 24117, 27366, 28764, 
    28717, 30049, 29820, 30528, 29469, 28895, 25077, 23017, 21454, 15869, 
    13499, 6805, 5902, -903, -3158, -9409, -13222, -17589, -21764, -21726, 
    -24850, -27552, -28953, -31058, -32346, -30347, -29571, -27865, -26515, 
    -23121, -20521, -15446, -12705, -9142, -4998, 228, 3392, 9709, 11238, 
    17249, 20576, 23229, 25684, 27022, 31302, 30129, 30932, 30225, 29693, 
    29286, 27028, 22658, 20360, 15594, 13092, 8813, 4421, -372, -5055, -7333, 
    -12577, -16821, -20211, -23083, -25527, -29305, -30013, -28775, -31362, 
    -29474, -29904, -27020, -26871, -23246, -19578, -16676, -12013, -7774, 
    -5066, 312, 5317, 9325, 13210, 16369, 20397, 24050, 25365, 27478, 29136, 
    30411, 31585, 30192, 30721, 27735, 27780, 25463, 19468, 17020, 13263, 
    7473, 4384, 1684, -5004, -8134, -11550, -16971, -19171, -21465, -26047, 
    -27825, -28172, -29911, -30833, -31525, -28273, -27478, -26512, -23228, 
    -20997, -17462, -13744, -9886, -5025, -1327, 2448, 7881, 10943, 15330, 
    20390, 23150, 24687, 28561, 27992, 29222, 29395, 31624, 29261, 29386, 
    27038, 23203, 21068, 16279, 15149, 8418, 5481, 346, -4492, -7437, -12977, 
    -15545, -18550, -22538, -25368, -27588, -28723, -29325, -30634, -30749, 
    -30182, -28889, -26643, -24367, -20935, -17922, -14526, -9555, -4973, 
    -456, 3316, 6093, 10916, 14413, 17777, 21577, 24394, 28495, 28936, 30091, 
    30870, 29190, 30285, 29269, 25716, 23464, 21008, 18551, 12949, 10231, 
    5196, 948, -3092, -5978, -12310, -14635, -19628, -22038, -25424, -25764, 
    -28514, -30431, -30830, -29883, -29171, -29267, -26358, -25550, -20014, 
    -18487, -14836, -11326, -6940, -1427, 4184, 6095, 10018, 14037, 19740, 
    21544, 24976, 28053, 29730, 29184, 31671, 31742, 31453, 29361, 28098, 
    24190, 22739, 18711, 14040, 10596, 5566, 2148, -3125, -6870, -9830, 
    -14030, -17591, -21978, -23377, -26230, -29356, -29812, -31235, -32318, 
    -29479, -28556, -27552, -24624, -22141, -19109, -13718, -9737, -5446, 
    -2305, 2615, 5196, 11278, 14581, 18586, 22609, 23460, 26987, 29646, 
    31420, 31397, 32050, 30330, 29940, 27919, 24716, 23662, 18420, 13910, 
    10021, 5837, 3780, -1202, -5560, -9704, -14555, -19772, -22058, -23832, 
    -26860, -28587, -29530, -31451, -30840, -30285, -28797, -26709, -24150, 
    -22178, -18939, -13687, -12072, -7723, -3763, 836, 4709, 9993, 15750, 
    18918, 21266, 25270, 25813, 27969, 29164, 30375, 32359, 31164, 30127, 
    27047, 24610, 22367, 19378, 15314, 11179, 8262, 4496, -1625, -5543, 
    -9841, -14088, -17783, -21304, -24285, -26733, -27642, -30501, -31420, 
    -31849, -31825, -28953, -28547, -25989, -23232, -20372, -14455, -13022, 
    -7763, -2940, 812, 6610, 10432, 13468, 17661, 21718, 24504, 27086, 29777, 
    30979, 31803, 32582, 29766, 27974, 28382, 25945, 23457, 20024, 15824, 
    11949, 7838, 2821, -1137, -5413, -9700, -13815, -16453, -20170, -22469, 
    -28011, -27456, -30223, -30461, -29531, -30342, -29930, -27114, -24421, 
    -21389, -20004, -14914, -12595, -7496, -3321, 824, 5866, 9030, 11879, 
    18601, 20880, 22601, 26497, 27918, 29617, 31746, 29628, 30962, 29771, 
    26336, 25356, 24375, 19467, 16298, 11553, 8792, 5485, -1356, -5830, 
    -8886, -13300, -16637, -21190, -22229, -26619, -28290, -28779, -30761, 
    -31053, -31012, -28434, -28190, -25011, -23987, -19459, -17572, -13104, 
    -7359, -3741, -709, 5539, 8191, 13457, 17271, 20126, 23180, 26803, 29204, 
    29809, 30019, 31836, 30567, 29701, 27924, 26992, 23132, 19058, 17177, 
    12344, 9471, 4167, -312, -3377, -8159, -13796, -17925, -20405, -22386, 
    -26762, -28053, -29490, -31546, -29755, -30237, -28797, -27463, -25113, 
    -23665, -21206, -15943, -12797, -9022, -5335, -1865, 4260, 8221, 12509, 
    16453, 20979, 22533, 25978, 27640, 28890, 30872, 30117, 29914, 27914, 
    28673, 25830, 23613, 19516, 18215, 13312, 10061, 4257, -32, -4320, -9008, 
    -14285, -16017, -20645, -23591, -26739, -26989, -30333, -31595, -29374, 
    -29561, -30014, -28062, -25926, -23430, -19002, -15505, -13543, -8869, 
    -3461, -178, 2609, 8509, 13493, 15941, 20344, 22933, 26304, 29642, 28058, 
    29584, 30838, 30473, 28649, 26904, 27423, 22891, 21515, 17687, 14780, 
    8184, 6457, 964, -3892, -7845, -11896, -14189, -20032, -22056, -26653, 
    -26970, -29453, -32176, -29878, -30595, -28845, -29439, -27568, -25287, 
    -19923, -18181, -13467, -9458, -5352, 18, 3180, 8195, 11887, 15386, 
    18836, 22147, 25433, 26308, 29540, 29664, 31846, 29905, 30104, 29754, 
    26367, 23333, 19910, 16973, 12901, 9524, 5395, 1032, -2973, -8219, 
    -12518, -15812, -20416, -21251, -24932, -27426, -29225, -30780, -31274, 
    -30459, -29205, -28377, -26572, -25179, -22174, -19002, -15634, -10105, 
    -5504, -786, 2422, 8323, 11515, 14768, 18903, 21887, 26443, 27367, 29366, 
    30420, 31048, 31261, 29371, 29583, 27008, 24782, 20833, 18803, 13081, 
    8853, 7205, 1933, -1953, -6272, -10789, -15396, -18785, -22729, -25058, 
    -27575, -29116, -28946, -32075, -31291, -30657, -28272, -27458, -23970, 
    -20616, -18767, -13861, -11527, -6249, -1688, 3319, 7661, 12243, 14322, 
    18608, 22186, 24055, 26652, 29113, 31518, 30613, 32233, 28841, 28447, 
    26775, 25963, 21354, 17251, 13783, 9399, 5781, 3200, -882, -5852, -11417, 
    -15411, -18618, -23247, -25282, -27191, -28788, -28905, -30198, -30832, 
    -29090, -29456, -25671, -23353, -22459, -17781, -14031, -9345, -5778, 
    -2409, 2372, 7755, 10765, 14026, 18483, 21105, 25364, 27300, 29672, 
    31252, 29036, 29501, 30427, 29078, 26202, 25416, 21708, 18346, 15113, 
    10674, 5218, 1845, -2079, -6888, -10138, -16366, -18379, -20163, -24376, 
    -27878, -27759, -28760, -30173, -29020, -29499, -29733, -27901, -24205, 
    -22673, -19790, -15078, -11368, -6080, -2842, 1321, 5841, 10664, 14515, 
    18225, 21726, 25379, 27645, 28393, 30130, 30199, 32272, 31290, 29239, 
    26829, 25816, 21481, 19369, 15245, 11321, 6757, 3248, -1546, -5942, 
    -10180, -15151, -18015, -21197, -24004, -25071, -27533, -29824, -31412, 
    -29253, -32070, -29284, -28188, -25411, -22608, -18901, -15692, -10673, 
    -7763, -3094, 910, 4756, 10562, 13643, 18694, 21185, 24823, 26006, 27435, 
    30108, 30570, 30660, 28759, 29215, 26647, 26160, 21148, 20723, 16084, 
    11522, 6923, 4350, -317, -4978, -10017, -13593, -16194, -19693, -23762, 
    -25855, -30292, -28894, -30551, -30414, -30398, -28275, -27309, -27067, 
    -21891, -18101, -15718, -13600, -7310, -2079, 1936, 4885, 9309, 14205, 
    17639, 20586, 24150, 26962, 29951, 29428, 31182, 31604, 30615, 29098, 
    28692, 25120, 21170, 19796, 14841, 10991, 8776, 3565, -728, -5102, -9142, 
    -11940, -17770, -18963, -24527, -26378, -28384, -30442, -30138, -29116, 
    -31583, -28856, -29275, -26399, -22500, -21025, -16073, -13780, -8418, 
    -4373, -24, 3377, 8728, 13695, 16556, 20812, 24827, 27719, 28004, 28671, 
    29704, 32085, 29897, 29467, 27749, 25852, 24505, 19916, 16500, 12338, 
    9353, 2434, 688, -4667, -8467, -14489, -16453, -20187, -24476, -26754, 
    -27324, -30132, -32220, -30177, -30155, -27922, -26695, -25825, -23569, 
    -20359, -17210, -13342, -8560, -6152, -931, 4547, 10046, 12996, 15429, 
    21768, 24311, 25327, 26961, 30443, 31435, 30752, 31711, 29641, 27687, 
    26732, 23078, 21324, 16642, 14220, 9946, 4855, 419, -5628, -9280, -12385, 
    -16841, -20510, -23392, -24995, -28469, -29947, -30507, -30400, -29130, 
    -29769, -29354, -25957, -24480, -21688, -18082, -11525, -9356, -4971, 
    -358, 2592, 9848, 12945, 14755, 21112, 24139, 25405, 28540, 28897, 30677, 
    29327, 30950, 31280, 27188, 27123, 22635, 21352, 18776, 13719, 10352, 
    6106, 1891, -4844, -8793, -11611, -16124, -19402, -23559, -25109, -27728, 
    -30438, -30212, -31979, -30469, -30126, -29165, -26850, -22601, -19242, 
    -17501, -13227, -9939, -4176, -2374, 4602, 9125, 10387, 15118, 20284, 
    21990, 25070, 28963, 29855, 30491, 29648, 30339, 29831, 28333, 24913, 
    22413, 19979, 18126, 14082, 10401, 4697, -249, -3353, -7842, -10922, 
    -15432, -17748, -23368, -26192, -26416, -29329, -29513, -31121, -29891, 
    -29807, -27785, -25886, -25103, -20723, -17976, -14729, -10524, -6140, 
    -1393, 2606, 6323, 11264, 16312, 18382, 22694, 24563, 28242, 29611, 
    28928, 32166, 30812, 28827, 27208, 27153, 25426, 20998, 17998, 14462, 
    11010, 5972, 582, -2542, -7413, -11357, -14162, -19323, -23076, -25640, 
    -27049, -28359, -30655, -30482, -29679, -29396, -29732, -25804, -24362, 
    -22094, -18333, -15136, -10629, -6009, -1522, 3385, 7370, 10153, 13998, 
    19178, 21540, 24773, 27359, 30202, 30032, 32012, 31082, 30354, 27333, 
    27183, 22978, 21036, 18427, 14734, 10847, 5785, 2353, -2717, -7585, 
    -10712, -16467, -19210, -21320, -24775, -25744, -28950, -30148, -30719, 
    -30583, -30275, -28222, -27726, -26301, -21698, -18496, -14748, -11670, 
    -7284, -3371, 3411, 6070, 10137, 13395, 18172, 22092, 24276, 26869, 
    28918, 31041, 32068, 30647, 30883, 29299, 27892, 23421, 21411, 17965, 
    13993, 12255, 6739, 2495, -2191, -6979, -10127, -14901, -17903, -21848, 
    -23315, -26463, -28373, -28906, -32225, -31989, -30294, -28420, -26577, 
    -24797, -21296, -18939, -13877, -12275, -6799, -3010, 2169, 6784, 11110, 
    13324, 18365, 22414, 23656, 25048, 28695, 30488, 30293, 30345, 30216, 
    29619, 25658, 24039, 22017, 18837, 14398, 11101, 6711, 3566, -2664, 
    -4619, -11486, -15370, -16522, -21304, -24026, -26615, -28052, -29244, 
    -29594, -30632, -29649, -28406, -26432, -25186, -23664, -18650, -16045, 
    -9901, -7418, -3054, 1374, 5784, 9240, 13075, 18282, 20248, 23527, 25244, 
    28602, 29962, 31819, 32433, 30216, 28830, 26811, 25217, 22493, 20002, 
    14802, 11451, 8290, 2889, -1507, -4229, -9411, -12024, -16351, -20802, 
    -24266, -26450, -28742, -30439, -29878, -31441, -29466, -27848, -29152, 
    -25470, -22937, -19444, -16140, -10729, -7860, -2883, 1771, 5196, 9553, 
    12979, 17052, 21599, 23994, 27209, 27434, 29579, 31417, 30452, 29182, 
    29386, 26694, 26640, 22903, 19389, 15575, 12514, 6331, 5009, -56, -5415, 
    -9074, -13193, -16956, -20504, -23566, -25337, -28162, -30592, -30543, 
    -29744, -30880, -29389, -29324, -25230, -22616, -19068, -16245, -12812, 
    -6637, -2943, 1388, 5041, 8885, 14489, 17018, 21603, 23636, 25726, 28768, 
    28791, 30458, 29723, 31271, 29158, 29054, 26866, 21987, 19571, 17092, 
    12613, 8091, 4520, -746, -3104, -7511, -13347, -16704, -20529, -23909, 
    -26313, -28795, -28984, -30911, -30856, -28759, -28849, -29124, -27256, 
    -22998, -20371, -16692, -13057, -8418, -3672, -859, 4535, 7499, 11969, 
    16167, 19930, 23834, 24275, 28047, 30575, 30063, 30406, 32132, 30030, 
    28034, 26331, 24660, 21289, 15805, 12646, 8140, 3399, 1098, -3009, -8509, 
    -12237, -17679, -20385, -22743, -25549, -28720, -28915, -30519, -31308, 
    -29245, -29234, -28400, -26053, -22662, -21505, -17332, -12733, -9500, 
    -4973, -128, 4838, 8552, 11270, 15624, 20112, 22900, 26869, 28320, 29622, 
    31543, 31467, 31235, 28491, 28505, 25958, 23729, 20356, 17318, 13269, 
    9468, 4512, -256, -2606, -8782, -13107, -17456, -20822, -23949, -25642, 
    -28448, -29366, -31833, -31639, -30849, -29981, -28856, -27914, -24361, 
    -22163, -17324, -13735, -9016, -4172, -2438, 3533, 7358, 10828, 14967, 
    20637, 23311, 25475, 28302, 29172, 30529, 32212, 30128, 29077, 29035, 
    25302, 23910, 21586, 17873, 13502, 9097, 6593, 1808, -1756, -7997, 
    -11690, -14985, -18442, -22100, -24121, -28540, -28812, -29846, -30251, 
    -31297, -28338, -27046, -26822, -23882, -20590, -17376, -13440, -9001, 
    -6145, -1161, 2246, 7382, 11468, 14883, 19161, 22925, 25857, 27414, 
    30148, 30034, 31387, 32168, 30109, 27676, 27947, 24531, 23084, 18403, 
    14689, 10426, 4568, 1950, -2134, -7596, -10941, -16952, -20165, -22187, 
    -25758, -27714, -29519, -31319, -29401, -29033, -28999, -29240, -27423, 
    -24666, -22746, -18581, -15531, -11020, -6738, -2571, 4039, 6583, 10174, 
    15398, 18164, 21246, 24326, 26481, 29540, 29726, 29693, 30047, 30332, 
    27250, 27035, 23127, 21413, 18640, 14263, 9825, 6865, 785, -3269, -6216, 
    -11015, -15471, -19377, -20949, -24280, -27258, -28723, -29801, -31978, 
    -29103, -30913, -29846, -27721, -23779, -22778, -17828, -14146, -11359, 
    -5795, -3302, 2555, 6604, 10831, 13658, 18465, 21329, 24817, 27915, 
    29953, 30259, 29849, 29842, 29230, 30455, 27184, 26335, 22129, 18552, 
    14567, 11902, 5627, 2897, -1011, -5345, -11367, -14856, -19146, -21746, 
    -23411, -26220, -29724, -31672, -30966, -32017, -30126, -29197, -27501, 
    -23592, -20938, -19292, -13478, -12253, -7089, -1325, 1787, 5925, 9259, 
    12869, 18091, 21464, 24393, 27676, 29242, 31271, 30365, 29795, 28811, 
    28635, 27086, 25297, 22596, 19238, 15646, 11221, 6653, 2713, -2025, 
    -5701, -9472, -14172, -19060, -22698, -23458, -26798, -30165, -28238, 
    -30520, -30875, -30879, -30428, -27513, -24569, -22526, -19145, -16763, 
    -10256, -7065, -3515, 2279, 6132, 8828, 13261, 18419, 21946, 23524, 
    28076, 29079, 30869, 30466, 31713, 31000, 28958, 26863, 26970, 21546, 
    19514, 15310, 10488, 6403, 2908, -1869, -6076, -9722, -13598, -18033, 
    -20864, -23887, -24664, -30187, -30541, -30565, -30378, -29975, -29083, 
    -27230, -24315, -23730, -19961, -15764, -12338, -7411, -2630, 2442, 6042, 
    8386, 12286, 18187, 19673, 24222, 26816, 27512, 30422, 30654, 32403, 
    28732, 28602, 27167, 24677, 24251, 19728, 16514, 11032, 7379, 3198, -440, 
    -6534, -7575, -13506, -15712, -20779, -24475, -26993, -29468, -30757, 
    -29415, -29364, -30814, -28465, -28883, -24927, -23205, -20300, -15715, 
    -11620, -6704, -3346, -656, 5055, 9144, 14056, 18661, 19768, 23790, 
    26898, 28498, 29194, 28907, 30195, 31535, 29300, 27816, 26479, 23893, 
    19298, 14786, 12514, 9699, 4160, -462, -4332, -7202, -12068, -16275, 
    -20185, -23037, -26271, -28587, -28241, -30724, -31071, -30662, -28262, 
    -28408, -25255, -24429, -20343, -16044, -14151, -8118, -4081, -1246, 
    4085, 7455, 12999, 16669, 19501, 23655, 26616, 29614, 30109, 31923, 
    30967, 32325, 29996, 27854, 26722, 23268, 19585, 16292, 12146, 9951, 
    2838, 1343, -3921, -8545, -13080, -17185, -19534, -23379, -25110, -27011, 
    -28851, -29574, -30543, -29820, -29206, -28240, -27270, -22997, -20243, 
    -16879, -13697, -8171, -4573, -581, 4061, 8503, 12060, 16594, 20866, 
    22153, 24620, 28660, 27571, 30896, 32307, 30074, 30693, 29031, 25655, 
    22947, 20433, 16529, 13157, 9295, 5319, 1225, -4116, -8448, -10948, 
    -15911, -20336, -22337, -24649, -27389, -31131, -30124, -29737, -31544, 
    -30445, -29222, -27359, -23545, -20895, -18212, -13627, -9284, -4221, 
    -1751, 3919, 8394, 11214, 16577, 19374, 22378, 26417, 27898, 29764, 
    31246, 30509, 30611, 29975, 27138, 25258, 22573, 20135, 17409, 13328, 
    9401, 5791, 117, -3243, -8111, -11139, -15209, -18174, -22578, -25066, 
    -28675, -30503, -30724, -31742, -30797, -31304, -28830, -25608, -24129, 
    -19364, -17669, -12410, -9499, -4810, -1108, 3983, 8812, 11081, 15663, 
    19545, 23994, 25148, 26087, 27998, 29358, 30989, 29460, 29821, 28114, 
    26526, 23615, 20726, 16639, 14423, 9863, 5936, 1299, -2838, -7442, 
    -12242, -15257, -17544, -22571, -24676, -27510, -29752, -28934, -31585, 
    -30684, -31549, -29599, -27787, -24416, -20355, -18425, -14816, -12123, 
    -5938, -3492, 2986, 7868, 12148, 14593, 16892, 22342, 24608, 27560, 
    29695, 31615, 30972, 29147, 30215, 28682, 26270, 23842, 21141, 18003, 
    15570, 8988, 6628, 1728, -4034, -7632, -11855, -14074, -18080, -22575, 
    -23350, -27865, -28619, -30933, -30867, -32187, -30241, -28598, -26445, 
    -24622, -20944, -18212, -16416, -10585, -4816, -1019, 2398, 5995, 11557, 
    16120, 18275, 22619, 24879, 25525, 28721, 30179, 30876, 30796, 31041, 
    29556, 27017, 24947, 21535, 17845, 15905, 9965, 6913, 2311, -2513, -6476, 
    -9055, -14242, -18702, -21409, -24527, -27846, -29447, -30289, -29533, 
    -32135, -28925, -28776, -27198, -24958, -21076, -18223, -15785, -10718, 
    -8218, -2897, 569, 7488, 11084, 15135, 17087, 20488, 23004, 25728, 29621, 
    30759, 31590, 31024, 31560, 28700, 27025, 26041, 21298, 18241, 16710, 
    10958, 8332, 2156, -1425, -5825, -9301, -14575, -16476, -21477, -24076, 
    -28357, -27739, -30007, -31760, -31387, -31438, -29410, -26903, -25560, 
    -22889, -18909, -15513, -12696, -7993, -3510, 1887, 6009, 11023, 13555, 
    18457, 21137, 22908, 26825, 28626, 29369, 31276, 30050, 29383, 29673, 
    27261, 26428, 22414, 18351, 15282, 10309, 7110, 2043, -1477, -5926, 
    -10390, -13924, -17564, -20681, -22968, -24776, -28490, -30058, -28988, 
    -29903, -28644, -28698, -27317, -26888, -22725, -18210, -15927, -10971, 
    -7591, -3484, 236, 4574, 9403, 13354, 17359, 20875, 23442, 27520, 27221, 
    29405, 31384, 31519, 30635, 28104, 28213, 23962, 22606, 20797, 15836, 
    11204, 9166, 3538, 724, -4123, -10278, -13539, -17613, -20349, -22961, 
    -24359, -28006, -29006, -30101, -30069, -30322, -28793, -27848, -24795, 
    -23093, -19964, -15151, -14104, -8253, -4035, 801, 5913, 10449, 13002, 
    17017, 21292, 23449, 25424, 27713, 29096, 30548, 32137, 30467, 28756, 
    28137, 24601, 21610, 20085, 16569, 12297, 7724, 5652, 243, -3779, -7609, 
    -14071, -17577, -20072, -22745, -27230, -27317, -29993, -29872, -30786, 
    -29474, -29652, -28520, -25518, -23723, -19516, -17396, -12630, -7366, 
    -5653, 594, 4297, 9234, 13110, 15741, 21580, 22439, 27080, 28336, 29824, 
    29633, 30247, 30029, 31048, 26659, 26211, 23076, 19689, 15700, 13356, 
    9003, 4931, 35, -4239, -8566, -13061, -16728, -18833, -22374, -27255, 
    -28573, -29753, -30412, -29830, -29354, -29185, -27577, -26164, -22822, 
    -20882, -16502, -13478, -8949, -3438, -417, 4065, 6932, 11919, 16613, 
    20045, 22729, 26437, 27575, 28446, 30478, 30033, 31554, 29602, 27882, 
    25197, 24312, 19480, 17000, 14618, 8874, 4762, -505, -2925, -6992, 
    -12655, -15848, -18577, -22329, -25105, -28045, -29446, -30016, -30571, 
    -30148, -29767, -29326, -26775, -24660, -21369, -16863, -14626, -9372, 
    -4250, -337, 2693, 8110, 11907, 17214, 19061, 21390, 25560, 26070, 28534, 
    30259, 31641, 29083, 29869, 29416, 26539, 23048, 20193, 17372, 13712, 
    9795, 4753, 1929, -3789, -7763, -10285, -15105, -18553, -21140, -26226, 
    -27107, -28525, -30025, -29757, -29749, -29644, -29097, -27350, -24295, 
    -19998, -17928, -13296, -8806, -5513, -709, 2545, 7797, 12347, 16406, 
    17842, 23066, 23774, 28019, 27817, 30926, 30522, 31749, 30234, 28400, 
    26135, 25648, 21543, 17236, 13742, 10098, 7128, 2136, -2880, -5934, 
    -11223, -14325, -19843, -23208, -25706, -28148, -30724, -30502, -31031, 
    -30846, -30382, -29820, -27266, -23915, -20600, -16683, -14601, -9584, 
    -5579, -754, 2676, 7239, 11093, 14751, 18362, 21231, 25768, 26557, 30403, 
    28701, 29895, 30191, 28889, 28984, 25699, 23739, 21832, 18791, 15345, 
    10242, 7088, 2621, -3592, -5250, -10535, -15715, -18743, -21834, -24714, 
    -27086, -29167, -30264, -29816, -31006, -31217, -27983, -25221, -24360, 
    -21758, -18370, -15462, -9192, -6805, -1770, 1822, 5823, 9732, 14484, 
    19101, 21701, 23932, 27527, 29375, 30322, 31356, 30543, 30220, 27967, 
    27728, 24784, 20927, 17958, 14108, 10838, 6004, 2141, -1265, -6050, 
    -10494, -15413, -18083, -21624, -24107, -25811, -28884, -31310, -31669, 
    -30747, -31646, -29212, -27404, -24943, -22824, -20522, -14230, -11247, 
    -7475, -2342, 2866, 6143, 8583, 15079, 18050, 20972, 24899, 28050, 29688, 
    29900, 30824, 31524, 29352, 29060, 26109, 25786, 20820, 19135, 14965, 
    12103, 8578, 3195, -1345, -5307, -11277, -14941, -17701, -22501, -24367, 
    -25654, -27059, -30116, -30382, -30412, -30620, -27442, -27012, -25673, 
    -20678, -18814, -14996, -11697, -7783, -1760, 3174, 6915, 8950, 12239, 
    19092, 20994, 25110, 27651, 27851, 30032, 31478, 30246, 29209, 27557, 
    27333, 25397, 21835, 18413, 15024, 10917, 5907, 3467, -1077, -4933, 
    -9904, -13723, -17018, -19747, -24047, -25265, -26798, -30804, -31179, 
    -31438, -30112, -29237, -28967, -24141, -22524, -19274, -16815, -12719, 
    -8549, -3975, 33, 5104, 9059, 13887, 16535, 20138, 22774, 25305, 28025, 
    29342, 30975, 31390, 31864, 29473, 28452, 25827, 24141, 19301, 15076, 
    10963, 6669, 4286, -854, -5026, -9410, -11811, -16195, -20080, -22630, 
    -26719, -28066, -29638, -31742, -30328, -31402, -30048, -26506, -24554, 
    -24196, -19855, -15097, -11816, -8469, -4520, 1404, 5358, 7308, 12908, 
    16083, 19210, 23534, 25707, 26559, 29017, 29533, 30641, 31308, 29388, 
    27613, 26454, 22976, 20787, 15032, 12979, 7549, 4993, -493, -5370, -9037, 
    -13076, -17740, -21301, -23835, -26590, -26885, -31100, -30841, -30594, 
    -29897, -29789, -28805, -25884, -23933, -19719, -17070, -12819, -7686, 
    -5115, 1228, 5631, 8898, 13821, 16438, 19243, 24276, 25614, 27126, 29095, 
    31715, 30678, 31034, 28623, 28265, 24782, 22823, 20451, 16691, 14216, 
    7889, 4598, 105, -5485, -8547, -13356, -16972, -19620, -21954, -26899, 
    -28614, -29476, -29736, -29939, -29867, -29489, -28827, -26041, -23023, 
    -19275, -18880, -14009, -7951, -3542, 875, 3705, 8644, 12340, 17656, 
    20700, 23642, 24988, 26219, 28199, 30215, 31412, 31958, 29617, 27316, 
    26577, 23864, 20973, 18215, 13252, 8320, 4891, 1780, -3205, -9099, 
    -12407, -16272, -19425, -23634, -25231, -26747, -29793, -30150, -31218, 
    -30538, -28424, -28044, -26524, -23065, -20719, -16186, -14240, -9396, 
    -5320, 956, 3194, 8326, 13291, 15366, 20287, 22353, 25963, 27328, 28578, 
    31942, 31392, 31520, 29789, 30039, 26394, 23530, 20619, 17862, 14329, 
    8881, 5296, 572, -3484, -6877, -12733, -14561, -18258, -21561, -24716, 
    -26873, -28430, -30798, -30594, -30128, -29508, -28567, -25922, -23699, 
    -21271, -17223, -13722, -9727, -4814, 438, 3568, 8243, 11143, 15933, 
    18908, 23037, 25529, 27399, 29019, 29183, 30682, 30088, 30502, 29506, 
    26478, 25313, 20717, 19152, 13695, 10559, 5004, 1179, -2394, -8542, 
    -11122, -14753, -19500, -21106, -25105, -26449, -29193, -30220, -31426, 
    -30399, -31555, -27738, -27480, -24719, -20512, -17450, -13328, -11673, 
    -5698, -857, 1296, 8026, 10851, 14164, 17511, 23757, 25185, 26146, 28933, 
    30521, 31300, 31017, 29957, 30211, 26035, 23780, 21011, 18069, 14617, 
    10505, 6586, 2696, -2728, -8334, -12064, -16156, -18323, -22769, -25963, 
    -26142, -28796, -30111, -29491, -31963, -31763, -28736, -25792, -24783, 
    -20421, -17449, -14399, -11502, -6890, -2175, 2205, 6951, 11288, 15260, 
    18235, 20745, 24595, 27100, 30013, 31048, 31339, 30540, 29224, 28482, 
    27496, 24091, 20328, 18938, 14710, 10370, 5492, 3297, -925, -6456, 
    -10538, -15116, -19229, -20625, -24528, -28045, -28066, -29410, -31741, 
    -32014, -28674, -28364, -26999, -24495, -22038, -17999, -15153, -11329, 
    -6495, -2248, 303, 5717, 9575, 15458, 17334, 22330, 24444, 26512, 27682, 
    30647, 30266, 32405, 30018, 29310, 26760, 26031, 22618, 18693, 16098, 
    12492, 8222, 2512, -1680, -6567, -10290, -13933, -17149, -22680, -23780, 
    -26614, -28116, -30545, -30845, -30336, -29507, -28619, -28680, -24144, 
    -22574, -19505, -15331, -10537, -8168, -4060, 790, 5806, 8813, 13271, 
    17027, 21571, 22998, 25084, 27320, 30430, 31798, 30953, 31974, 29669, 
    28202, 25067, 23054, 19846, 15634, 11714, 7268, 2998, -1976, -4042, 
    -9529, -12769, -17881, -19191, -23488, -27303, -28921, -30610, -30722, 
    -31880, -30761, -29345, -27425, -23866, -22759, -19987, -15531, -13234, 
    -8533, -4580, 1820, 4433, 9767, 14432, 17446, 20862, 23832, 27562, 28926, 
    30622, 30725, 30627, 31383, 30496, 28123, 26509, 22809, 19620, 16052, 
    11979, 8028, 2105, -833, -5825, -8520, -13705, -16292, -21477, -23427, 
    -26808, -28401, -28573, -31802, -32382, -30423, -29115, -28845, -26247, 
    -22992, -19367, -16999, -12870, -6435, -4404, -945, 4604, 7919, 13023, 
    15849, 21068, 23637, 24353, 26817, 29919, 30374, 31959, 29173, 28742, 
    26826, 26147, 21964, 19984, 15214, 13291, 8599, 4348, 154, -4114, -9855, 
    -11666, -17728, -21500, -23168, -26836, -27803, -29092, -32250, -31627, 
    -30914, -28567, -28902, -25797, -21934, -20376, -16088, -12331, -8851, 
    -4268, 1409, 5219, 9443, 12914, 17022, 19919, 22860, 25114, 28294, 28222, 
    30399, 30675, 30615, 28391, 28602, 25404, 21648, 19725, 16276, 11779, 
    10173, 4236, -307, -2999, -7590, -13066, -15226, -19984, -24313, -25043, 
    -27869, -29325, -29737, -31683, -30880, -30315, -28787, -26126, -23352, 
    -22161, -18648, -13410, -8068, -4018, -326, 4315, 7848, 13771, 16002, 
    19598, 24206, 25804, 27111, 28910, 29659, 31857, 30945, 29596, 29514, 
    26537, 23752, 21550, 17926, 14852, 9470, 3593, 1112, -4789, -7913, 
    -12150, -15800, -20015, -23508, -25893, -27418, -29529, -29491, -31716, 
    -31071, -29655, -28876, -26496, -22075, -20192, -17942, -14541, -9926, 
    -5910, 716, 3744, 6764, 10139, 15257, 20273, 22879, 25753, 28955, 28956, 
    30550, 30580, 29650, 28998, 28045, 27376, 24321, 21249, 17736, 15026, 
    10097, 7022, 2607, -4595, -7590, -10618, -14734, -19190, -23396, -24778, 
    -28246, -28622, -31470, -31084, -30984, -29063, -27091, -26376, -25426, 
    -20294, -17796, -12927, -10064, -6783, -978, 3682, 7259, 13396, 16152, 
    18947, 21582, 26777, 27811, 27982, 31173, 30957, 30673, 29286, 27493, 
    27226, 23961, 19658, 16982, 15755, 10135, 7151, 582, -2879, -7846, 
    -12422, -15059, -19748, -22730, -25700, -26922, -27997, -31624, -30946, 
    -29874, -29846, -27439, -26573, -22640, -22055, -17323, -14885, -11428, 
    -6237, -1743, 2439, 6351, 11012, 15743, 19503, 21743, 24007, 28529, 
    29071, 28702, 31611, 30447, 28807, 28136, 26466, 24138, 20563, 19122, 
    14012, 10562, 6348, 309, -2958, -5428, -9378, -14485, -17806, -22468, 
    -24405, -28435, -28031, -31411, -30554, -30214, -30140, -29614, -26966, 
    -24773, -22131, -19475, -13689, -11229, -7515, -667, 1656, 6658, 10837, 
    14739, 18919, 22005, 25420, 28056, 27423, 30018, 32090, 30750, 30169, 
    30602, 27584, 24959, 22261, 18117, 15432, 11599, 6821, 2754, -1201, 
    -7464, -11927, -14192, -18338, -20734, -25097, -27281, -28995, -30316, 
    -29847, -29949, -31140, -28796, -28628, -25367, -21959, -20649, -14497, 
    -11658, -7246, -2326, 1266, 6168, 11053, 13345, 18300, 20123, 24201, 
    27316, 27684, 30781, 30991, 31589, 30824, 29006, 26035, 24388, 22259, 
    19254, 15925, 10454, 8028, 2593, -1039, -6006, -10451, -12550, -17621, 
    -19897, -24546, -25986, -28545, -30504, -30588, -30820, -30227, -29552, 
    -26685, -23848, -22335, -20191, -17033, -11679, -7011, -2482, 1765, 4987, 
    8513, 12410, 17822, 20207, 23125, 25070, 29679, 30922, 31373, 31410, 
    30687, 28898, 27799, 24764, 21481, 18715, 15837, 12217, 7484, 3225, -280, 
    -5521, -10885, -12951, -17232, -20554, -23933, -24935, -29411, -30323, 
    -30210, -31590, -32061, -29107, -27027, -24082, -22366, -20705, -16245, 
    -12906, -7937, -3442, 2094, 3837, 8533, 14128, 17079, 20047, 23457, 
    24924, 27282, 30231, 30156, 30700, 29525, 27771, 29534, 25226, 22149, 
    19541, 16140, 13057, 6904, 2150, -240, -4239, -10613, -12676, -17186, 
    -19860, -23668, -26313, -28162, -27973, -29769, -29562, -31019, -28338, 
    -28484, -25697, -22788, -19093, -17042, -12357, -7694, -4630, 938, 4012, 
    8930, 12512, 16842, 21265, 25015, 24356, 28164, 29278, 30340, 31204, 
    29720, 28137, 27406, 25302, 23253, 19947, 16085, 14013, 8154, 5018, 150, 
    -5124, -9791, -11682, -17306, -20096, -22581, -24923, -27746, -29583, 
    -30700, -30331, -31043, -29617, -28822, -25576, -23958, -19488, -16484, 
    -13189, -7713, -3350, -532, 4899, 8851, 14470, 16462, 19560, 23839, 
    24619, 28365, 27917, 31360, 30783, 30755, 28736, 27366, 26097, 23292, 
    20553, 18127, 12938, 8709, 6145, 50, -4016, -9590, -14103, -17151, 
    -20193, -23437, -24736, -27226, -30548, -30127, -30828, -30976, -29332, 
    -27345, -25684, -24309, -21387, -17558, -12602, -9224, -5783, -282, 4912, 
    9331, 11849, 16639, 19713, 22931, 24638, 27184, 31066, 30619, 29439, 
    29036, 30812, 27730, 25125, 22539, 19483, 18777, 13441, 10234, 5475, 
    1661, -5470, -8939, -10817, -16432, -19436, -23391, -24862, -29466, 
    -28442, -30265, -32006, -29841, -30325, -27973, -25814, -23202, -19945, 
    -18164, -13537, -9776, -5387, -1418, 1920, 7534, 11247, 17763, 19034, 
    23121, 24106, 27993, 30686, 30373, 30973, 28909, 30281, 28491, 26237, 
    24818, 20580, 16448, 13912, 9182, 5616, 1036, -4092, -7632, -13006, 
    -15895, -17741, -22401, -25412, -27940, -30603, -28867, -30611, -30654, 
    -29547, -29210, -26563, -24237, -22293, -18086, -13556, -9966, -6531, 
    -1165, 2937, 6069, 12843, 15894, 17511, 23130, 26121, 28827, 28086, 
    30513, 30545, 31811, 30818, 28478, 25719, 23251, 19752, 16881, 13544, 
    10234, 6452, 1789, -1356, -7931, -12359, -16777, -18380, -22439, -26103, 
    -29014, -29157, -29593, -30893, -31102, -29516, -28197, -26933, -25470, 
    -21597, -18681, -13624, -10931, -5821, -1731, 2191, 8204, 10108, 13747, 
    17773, 21108, 25722, 28054, 28525, 30585, 30910, 30736, 31167, 27859, 
    27078, 24373, 21941, 18634, 13993, 12039, 7043, 1068, -1508, -6972, 
    -9791, -14879, -17582, -21331, -25313, -26107, -28994, -29548, -31546, 
    -30287, -28894, -29136, -26329, -25651, -22114, -17198, -15728, -12332, 
    -6962, -2214, 1496, 4818, 10402, 15678, 18715, 23455, 25145, 27607, 
    29521, 31327, 30953, 29528, 29477, 30167, 26163, 25138, 20660, 19486, 
    16653, 11911, 7036, 4213, -2142, -5189, -11597, -14595, -17927, -22642, 
    -25482, -26833, -29599, -30624, -30596, -30094, -31032, -28883, -27037, 
    -25117, -21997, -19114, -15158, -10815, -6967, -2663, 987, 5582, 10406, 
    14396, 16441, 22057, 25277, 26018, 30023, 29881, 31233, 30550, 31028, 
    28278, 26925, 24412, 21758, 20387, 15582, 11969, 7584, 3932, -805, -5507, 
    -10550, -14256, -16998, -20791, -23445, -26194, -28738, -29940, -28853, 
    -31240, -31632, -30231, -27450, -25234, -23792, -19817, -16571, -12574, 
    -8100, -2767, 2935, 5501, 9908, 14112, 18289, 19634, 24392, 26507, 29402, 
    30076, 29314, 29668, 30208, 30728, 27509, 26205, 22007, 19236, 15165, 
    11209, 7913, 1765, -2092, -5253, -10239, -13339, -15897, -21608, -24553, 
    -26919, -28582, -30228, -29956, -31726, -30197, -28478, -27483, -24434, 
    -22083, -19855, -15583, -13353, -6994, -4963, -426, 5403, 9579, 12402, 
    17544, 19616, 22241, 27096, 27884, 30843, 30173, 30164, 30868, 29236, 
    27262, 24932, 24098, 19682, 16251, 12612, 7208, 3783, 51, -4088, -9083, 
    -14343, -16651, -20654, -24269, -27235, -26759, -31247, -31200, -29691, 
    -30336, -29565, -28597, -26391, -22729, -21195, -15819, -11967, -9506, 
    -4382, -713, 4721, 8257, 12675, 16203, 21343, 23649, 25796, 26514, 29692, 
    28905, 30922, 29278, 29873, 27419, 25153, 22040, 20042, 17292, 12298, 
    9919, 4134, 656, -4675, -8147, -13471, -18103, -18925, -23267, -24684, 
    -27330, -29454, -30352, -30612, -30808, -27902, -28520, -25381, -21790, 
    -20117, -17293, -12667, -9148, -4564, -162, 5465, 9454, 12815, 16201, 
    18701, 24130, 25285, 26616, 29584, 31815, 31594, 29633, 29333, 27408, 
    25881, 22968, 21137, 16993, 11499, 9187, 3112, 447, -4089, -7792, -11247, 
    -16211, -19620, -23590, -24300, -28941, -29856, -31079, -29751, -30674, 
    -31299, -28067, -27094, -23770, -21956, -16950, -12427, -10703, -4524, 
    -14, 4030, 9903, 12811, 15968, 19624, 22240, 27409, 28778, 27838, 30365, 
    31466, 29906, 29589, 28446, 25739, 23770, 20066, 16442, 14448, 10624, 
    5284, -1240, -5158, -8684, -11958, -16483, -19566, -21422, -23964, 
    -28988, -29140, -29365, -30038, -31053, -30050, -26844, -25227, -25409, 
    -21338, -17444, -13978, -9608, -5695, -1045, 3900, 7029, 12140, 16186, 
    20420, 21713, 25229, 27468, 29818, 31030, 31718, 30553, 30662, 28891, 
    27668, 24175, 20953, 16880, 14133, 8921, 5474, -443, -3033, -7477, 
    -11916, -13858, -18614, -21690, -25492, -28279, -28505, -29590, -31321, 
    -31501, -28687, -29102, -27177, -23238, -21794, -18928, -12144, -8769, 
    -5799, -699, 2626, 5959, 10582, 15409, 20423, 23399, 25704, 26524, 29075, 
    30217, 29430, 31078, 28780, 28794, 27563, 23785, 19978, 18930, 14465, 
    10667, 5356, 1426, -3330, -8509, -11522, -13891, -17855, -22088, -24858, 
    -28414, -27489, -30019, -29796, -30802, -31550, -28730, -27710, -23602, 
    -22806, -19110, -15615, -10596, -6786, -2360, 1594, 6603, 10485, 14846, 
    18672, 22547, 25221, 26976, 27830, 29522, 30531, 31902, 29556, 30107, 
    25795, 24452, 20994, 17439, 15056, 11919, 6243, 697, -1886, -6848, 
    -10345, -15537, -18347, -22833, -24252, -27696, -28034, -30114, -31542, 
    -30171, -30825, -27761, -27850, -23990, -22878, -17653, -12868, -9505, 
    -5755, -1795, 1741, 5786, 10757, 14928, 17867, 21152, 25460, 26017, 
    29773, 29139, 31168, 29983, 29602, 28622, 26533, 24412, 21513, 19186, 
    14940, 10339, 5285, 1837, -1939, -6805, -10429, -15831, -18351, -21376, 
    -25203, -27251, -29302, -28645, -31544, -31115, -30026, -28161, -27013, 
    -24014, -21176, -19156, -14365, -10193, -7768, -3239, 2664, 6679, 10111, 
    13323, 18137, 22313, 23518, 27165, 28473, 28528, 31634, 31364, 30698, 
    28741, 26907, 25524, 21518, 19247, 15810, 10950, 8651, 4052, -2622, 
    -5935, -10404, -15016, -18851, -21181, -24141, -25969, -26881, -30053, 
    -30148, -31814, -31049, -27979, -27321, -25216, -21573, -19088, -15540, 
    -11398, -6096, -2912, 1229, 4424, 9806, 14103, 18073, 22177, 22907, 
    26619, 28343, 28567, 30367, 32213, 30154, 28610, 27027, 24475, 22104, 
    17735, 15037, 12021, 7316, 2927, -1578, -6750, -9772, -12472, -15939, 
    -19634, -23964, -27601, -28001, -29921, -30539, -29868, -31410, -29661, 
    -26706, -25521, -23587, -19402, -14709, -11549, -7641, -4131, -574, 6257, 
    10084, 13145, 19198, 20836, 22708, 26320, 28196, 29307, 31066, 30411, 
    30112, 30038, 27891, 24890, 21644, 20470, 17661, 11808, 8723, 3271, 33, 
    -5588, -7864, -12834, -17030, -19739, -22809, -26951, -28390, -28128, 
    -30914, -31314, -29777, -29405, -28085, -25844, -21576, -21276, -15909, 
    -10975, -8332, -3758, 2003, 4480, 8053, 12161, 18250, 21038, 23712, 
    25171, 27643, 31165, 31847, 30873, 30816, 28485, 26825, 25614, 23167, 
    19744, 16787, 12895, 9645, 4244, -212, -5295, -9104, -13160, -16716, 
    -20945, -24641, -25715, -28464, -30854, -30701, -30992, -30007, -30326, 
    -27609, -25518, -21911, -20309, -16670, -12695, -9810, -4373, 50, 5340, 
    8698, 12827, 16496, 18697, 22429, 25296, 29108, 29744, 31380, 30908, 
    31185, 29784, 28024, 26025, 23735, 21243, 18192, 14361, 9376, 3443, -343, 
    -5061, -9341, -11957, -15902, -20154, -23164, -25483, -28647, -29719, 
    -29522, -32281, -30143, -28887, -28677, -25991, -23706, -21628, -17665, 
    -12018, -9390, -5598, -1259, 4931, 8203, 12366, 16902, 20082, 22088, 
    26180, 27701, 29662, 30672, 32333, 30827, 29449, 29256, 26945, 22790, 
    21899, 17814, 13199, 8847, 4388, -458, -4355, -7899, -10935, -16125, 
    -19053, -23113, -25110, -27103, -30012, -30518, -30373, -29390, -30992, 
    -29237, -25267, -23363, -20495, -17276, -13825, -9946, -5581, -68, 3468, 
    7858, 12242, 16902, 19661, 23736, 26064, 27819, 30651, 30475, 29758, 
    29624, 30353, 27523, 27204, 22220, 20273, 17614, 14967, 9230, 4093, -2, 
    -3459, -8494, -11418, -14391, -20283, -23172, -26346, -27671, -30823, 
    -30553, -31027, -29729, -29674, -27051, -26479, -25420, -20327, -18334, 
    -13436, -8907, -4939, -2139, 3564, 8075, 12777, 14322, 20228, 22657, 
    24828, 26205, 28721, 32079, 31439, 30732, 28847, 28137, 25534, 24010, 
    22606, 17647, 14778, 10087, 5391, 624, -2537, -6998, -11210, -14023, 
    -18239, -22713, -26361, -28871, -28969, -30340, -30930, -30258, -29923, 
    -29330, -27463, -24750, -20129, -17837, -12924, -11049, -7286, -2309, 
    2142, 5785, 11163, 14735, 19494, 21818, 24422, 25639, 28506, 29861, 
    31051, 31415, 29525, 28017, 27817, 25459, 21138, 17327, 14756, 10885, 
    5494, 1841, -1202, -6918, -11703, -14623, -17597, -21209, -24337, -26970, 
    -29245, -29516, -29658, -29795, -29293, -27886, -26411, -24211, -21793, 
    -18524, -14600, -10691, -6646, -3362, 3288, 4960, 10636, 15017, 19507, 
    21498, 23001, 26747, 27918, 28620, 31448, 30910, 30360, 29636, 26616, 
    25575, 20542, 18206, 15727, 12056, 7353, 2283, -497, -6193, -9894, 
    -16134, -17302, -20128, -24680, -27342, -29889, -29953, -30443, -31890, 
    -30098, -27236, -26033, -25587, -22397, -17642, -14996, -11294, -8388, 
    -2365, 3374, 5276, 9753, 13632, 18116, 22028, 24092, 27116, 29514, 29307, 
    29069, 29999, 28741, 29162, 26908, 25139, 23068, 18438, 14264, 11669, 
    7222, 3507, -1484, -5877, -10352, -13655, -16467, -21384, -25160, -27121, 
    -27984, -29858, -29777, -30917, -30710, -28490, -28506, -24897, -22510, 
    -17539, -16800, -10567, -5959, -2713, 970, 5827, 10606, 14586, 17420, 
    20237, 23940, 27668, 28069, 29832, 30902, 30127, 30892, 29437, 28522, 
    26310, 22906, 20405, 14779, 11338, 7003, 2519, -439, -5675, -10413, 
    -14128, -16833, -20468, -24972, -27542, -27260, -30021, -30810, -31659, 
    -29005, -29270, -27024, -25675, -23302, -19294, -16037, -13269, -8615, 
    -3386, 452, 4476, 9048, 13421, 18144, 20935, 23591, 26924, 28735, 31217, 
    32080, 30069, 29720, 29108, 27564, 23950, 21438, 18381, 15879, 11915, 
    8621, 3285, -63, -3879, -9255, -12709, -17964, -19476, -23569, -25338, 
    -26982, -30810, -31991, -30544, -30185, -28023, -28906, -25535, -22236, 
    -18734, -14985, -11448, -9405, -4207, 1506, 4490, 9724, 13813, 17390, 
    20713, 23019, 26416, 27825, 29655, 31882, 29902, 30766, 28776, 27054, 
    27560, 22587, 20742, 17609, 12616, 7896, 4397, 186, -3607, -7663, -12352, 
    -16800, -19278, -23862, -26039, -28784, -29673, -29772, -30374, -29820, 
    -28787, -28693, -24602, -22821, -18514, -16147, -11823, -9986, -5762, 
    -187, 5137, 7553, 14511, 17597, 18471, 22550, 25897, 28052, 29454, 29791, 
    30582, 31029, 30831, 27657, 24433, 23781, 19161, 18486, 13499, 7367, 
    3786, -331, -3973, -8341, -12812, -15483, -19915, -22307, -26646, -28464, 
    -30788, -31541, -30297, -30402, -28976, -28343, -26649, -23489, -21244, 
    -16718, -13119, -9020, -4000, -1105, 3473, 7604, 11381, 15563, 19620, 
    23770, 25863, 28049, 30248, 30791, 31115, 30332, 29089, 27633, 27833, 
    23915, 19566, 17888, 13617, 9224, 4862, 1398, -3419, -8903, -11781, 
    -16050, -19557, -22802, -24053, -27691, -29904, -30151, -29858, -31201, 
    -29016, -28785, -27106, -24440, -21142, -17113, -14966, -8532, -6648, 
    -1813, 3388, 7562, 12524, 16227, 20365, 22207, 25673, 26938, 29259, 
    30757, 31055, 30545, 29015, 28130, 25566, 25023, 22023, 17953, 14487, 
    9654, 4684, 791, -1580, -7022, -10403, -15631, -19770, -23852, -25906, 
    -28689, -30801, -31419, -31595, -30246, -28885, -27769, -26853, -25251, 
    -21454, -16417, -15655, -11036, -5460, 16, 2828, 6914, 12128, 16860, 
    20659, 22824, 25085, 28411, 30833, 30488, 30590, 30448, 28623, 28294, 
    27183, 25657, 19618, 17210, 13365, 10222, 4967, 1187, -1645, -6068, 
    -11492, -15718, -17661, -21777, -25023, -27505, -29182, -29640, -32458, 
    -30690, -30924, -29880, -27022, -24936, -21270, -18012, -14227, -9383, 
    -7236, -1355, 3815, 7872, 12401, 14043, 17238, 21998, 25307, 26839, 
    30252, 31778, 30120, 29803, 29959, 29581, 27136, 25464, 22092, 19284, 
    15465, 9317, 7059, 1657, -3467, -5667, -12412, -16379, -19905, -20220, 
    -24818, -27158, -28130, -30221, -31271, -30166, -31526, -27872, -26262, 
    -24408, -22227, -18199, -15033, -12066, -5065, -2058, 2572, 6100, 11990, 
    14076, 19478, 20114, 23725, 27873, 28144, 29116, 29372, 31022, 30681, 
    27949, 27686, 23442, 22631, 17794, 14607, 10620, 6440, 1804, -1064, 
    -6375, -12050, -14852, -18360, -22680, -24413, -27972, -28816, -30049, 
    -30838, -30060, -30767, -29195, -28188, -25561, -22139, -18640, -15258, 
    -10719, -6450, -2509, 527, 6209, 9453, 13747, 18143, 21991, 23696, 25815, 
    28852, 30041, 31840, 30605, 30693, 28864, 26346, 25421, 22480, 19614, 
    16125, 11626, 8077, 2222, -1978, -5101, -10498, -14329, -18675, -21614, 
    -23661, -28100, -27501, -31380, -30820, -29735, -30874, -28588, -27944, 
    -24993, -20743, -17895, -14317, -10276, -7465, -4284, 1227, 5687, 10141, 
    15580, 17761, 21303, 24422, 27125, 28609, 30315, 31261, 29555, 30517, 
    28804, 28106, 25799, 23978, 19092, 14592, 13086, 6363, 2492, -475, -4629, 
    -11151, -13806, -16870, -21076, -22829, -26499, -28576, -30965, -30819, 
    -30937, -31285, -29749, -28403, -25720, -22053, -20950, -15976, -11059, 
    -8238, -3615, 950, 5539, 9271, 13458, 16059, 19478, 23945, 26815, 28489, 
    29431, 30640, 29674, 29185, 29292, 26068, 25720, 23101, 18403, 15761, 
    10452, 7285, 2596, 178, -4188, -9722, -12015, -17265, -19028, -22757, 
    -26360, -27000, -31015, -30064, -31053, -30048, -30556, -27710, -24093, 
    -23589, -20061, -17334, -12683, -7520, -4804, 190, 4894, 9487, 12753, 
    15936, 20785, 23586, 25174, 27437, 30086, 29692, 31346, 31359, 29085, 
    28253, 25487, 22889, 20213, 17207, 12059, 7368, 3850, -57, -4116, -8955, 
    -13776, -17800, -19298, -21639, -25453, -28140, -31235, -29517, -30429, 
    -31492, -30168, -28670, -24430, -23599, -20801, -17738, -12667, -9417, 
    -4934, -877, 2905, 6845, 13013, 15585, 21133, 22202, 26492, 28425, 29370, 
    31234, 30804, 30650, 29466, 27554, 26237, 23098, 19870, 17634, 12095, 
    9058, 5450, 129, -3227, -8622, -13530, -15324, -18739, -23918, -26360, 
    -29241, -31056, -30579, -30489, -31113, -28811, -27251, -24967, -24866, 
    -21937, -16532, -13275, -9226, -4404, 341, 4054, 7423, 11579, 15610, 
    19660, 23538, 25669, 28548, 28946, 29600, 30543, 29360, 29349, 27549, 
    25252, 24866, 20411, 17922, 11708, 10347, 6378, 1066, -4452, -7601, 
    -12394, -15224, -18211, -22493, -25846, -26627, -30407, -30402, -32307, 
    -30066, -30026, -26857, -25671, -23455, -21072, -17089, -13291, -8903, 
    -6212, -525, 3512, 6481, 12515, 15944, 20167, 23684, 25406, 26176, 29170, 
    29669, 29791, 30549, 29591, 28986, 26389, 23279, 21828, 17802, 14350, 
    9468, 6808, 1174, -3460, -6503, -12374, -16295, -18497, -22194, -24117, 
    -27287, -29034, -29348, -29859, -30711, -29776, -29742, -24897, -25157, 
    -20747, -17762, -13918, -11645, -6049, -1381, 3156, 6050, 11745, 16167, 
    20374, 21340, 25720, 27563, 28545, 30419, 32003, 31556, 31021, 29373, 
    26645, 22742, 21512, 17876, 14778, 11050, 5140, 1435, -3044, -8785, 
    -11053, -15524, -18647, -21009, -24893, -27918, -28249, -29206, -30960, 
    -30712, -29364, -28905, -26228, -23556, -21465, -16913, -13451, -11120, 
    -6203, -2094, 3719, 6734, 10869, 15343, 20139, 21792, 24624, 27738, 
    30487, 31315, 30472, 32564, 30012, 27900, 27555, 24661, 21980, 19208, 
    14816, 10387, 6228, 1578, -2713, -6840, -10404, -15288, -18700, -22879, 
    -26194, -27470, -29266, -29961, -30100, -29280, -29410, -29655, -28315, 
    -25206, -20982, -18407, -16091, -10349, -6598, -3684, 2335, 6821, 11024, 
    13306, 17515, 20941, 26105, 25889, 28224, 30451, 30402, 29164, 31062, 
    27963, 28568, 24374, 22572, 18540, 15284, 10295, 7724, 1606, -2385, 
    -5487, -10501, -13584, -18992, -19886, -23318, -26592, -30097, -30931, 
    -30354, -30004, -30140, -28876, -26874, -24783, -21898, -18196, -14003, 
    -9962, -6068, -2190, 3183, 6731, 10174, 13412, 17950, 21907, 24274, 
    26660, 30006, 29962, 31605, 31597, 31703, 29446, 27739, 23118, 22311, 
    18566, 15230, 12186, 7313, 2852, -2670, -7071, -9581, -14128, -18026, 
    -21580, -23945, -27544, -28751, -30451, -30795, -30583, -30211, -29767, 
    -26869, -25420, -22237, -20503, -16514, -10549, -7985, -2412, 2360, 5199, 
    9632, 15081, 17708, 21992, 23981, 25395, 27485, 29299, 30164, 31090, 
    30216, 28326, 27759, 25922, 22303, 20247, 16495, 10562, 7535, 2707, 
    -1774, -4825, -10382, -15617, -16635, -20645, -22912, -26855, -28870, 
    -29927, -29938, -32452, -29918, -29863, -26048, -24534, -22029, -19535, 
    -15663, -11627, -8889, -4991, 1464, 4707, 10356, 13628, 15986, 20514, 
    24009, 25948, 29670, 29683, 31248, 31735, 30932, 29378, 27884, 25416, 
    23734, 20443, 16143, 12280, 8453, 4409, -624, -5881, -9530, -13092, 
    -16826, -19296, -22186, -25907, -28357, -30599, -29679, -29547, -31000, 
    -28988, -28098, -25408, -22643, -18594, -16374, -13000, -8976, -3641, 
    -721, 4747, 8786, 13227, 16798, 20353, 25033, 24985, 28398, 30290, 30379, 
    31388, 29615, 29242, 27054, 25937, 23456, 18800, 15878, 12588, 7596, 
    3036, -744, -4230, -8730, -13423, -17201, -19256, -22160, -24571, -29859, 
    -30790, -31929, -30569, -31095, -29896, -29098, -25952, -22700, -20532, 
    -16572, -12755, -9468, -4267, 463, 4331, 7721, 14089, 14842, 21219, 
    23515, 24910, 29374, 29778, 31112, 31207, 29448, 30101, 28463, 24436, 
    22687, 20256, 15453, 13399, 7216, 4038, -648, -4681, -9006, -12384, 
    -16649, -19972, -23158, -26940, -28437, -29486, -29929, -31221, -30340, 
    -29689, -27745, -25418, -24190, -20625, -16959, -13506, -8544, -5714, 
    -1478, 2070, 7293, 12807, 15872, 20220, 22575, 24984, 28318, 29299, 
    31141, 31121, 31266, 29567, 28095, 25845, 23569, 21507, 17233, 13918, 
    9374, 4374, -498, -2636, -7324, -13050, -16576, -19265, -23538, -26212, 
    -26908, -28432, -31118, -31615, -28757, -29224, -28340, -27725, -23524, 
    -19373, -17646, -13550, -9384, -6219, -946, 3523, 7101, 13826, 15739, 
    19702, 21033, 25498, 27453, 29147, 31242, 30628, 31087, 29485, 28036, 
    26877, 23287, 20314, 18615, 14340, 10548, 6178, 506, -3201, -7347, 
    -11632, -15856, -18365, -22159, -24990, -26415, -28908, -29971, -30857, 
    -29931, -31347, -26735, -25850, -24468, -22186, -17230, -14111, -9292, 
    -4584, -2122, 2837, 7871, 11310, 13975, 19070, 21364, 25685, 28150, 
    28856, 30134, 29119, 30759, 30675, 27933, 26551, 23252, 22391, 17583, 
    15216, 11317, 4703, 458, -1920, -7316, -10993, -14027, -19635, -23301, 
    -25040, -27205, -28978, -29915, -29882, -29637, -29849, -29805, -25543, 
    -24329, -22054, -18192, -13403, -10675, -5663, -2527, 2716, 6795, 9393, 
    15182, 19732, 21640, 25001, 27012, 28715, 28544, 31542, 30607, 31067, 
    27610, 26512, 24205, 22522, 17745, 14354, 9987, 6843, 2213, -2919, -5935, 
    -9410, -14980, -18980, -22602, -25244, -26002, -28999, -30745, -30905, 
    -30230, -30081, -28781, -26792, -23965, -21584, -17214, -14834, -9180, 
    -6932, -2278, 906, 7920, 10812, 14426, 19813, 20591, 25880, 26991, 28890, 
    30892, 30254, 31359, 31108, 29226, 26974, 24708, 22129, 19319, 14923, 
    11299, 6453, 963, -2550, -6790, -11184, -15597, -18149, -20721, -23962, 
    -27469, -29846, -30114, -29548, -30231, -29177, -27471, -27158, -24676, 
    -20518, -19323, -16233, -9532, -6923, -4142, 1449, 6817, 8984, 13221, 
    18130, 22168, 24325, 26672, 29975, 30881, 31092, 31646, 30939, 29192, 
    26072, 24989, 23034, 19313, 13620, 11310, 7722, 2409, -2680, -5762, 
    -10529, -14283, -16165, -21919, -25763, -27002, -29684, -29416, -30823, 
    -31919, -29827, -28216, -27512, -25573, -21279, -19464, -15119, -12705, 
    -8297, -2403, 174, 5827, 8725, 13646, 17662, 20196, 25297, 26522, 29180, 
    29693, 30375, 30888, 30946, 29072, 28433, 26406, 22682, 19024, 15570, 
    12913, 7288, 3526, -1139, -6126, -10922, -12244, -18709, -21482, -23366, 
    -27064, -27036, -30437, -30570, -31880, -31220, -28046, -28574, -25323, 
    -23269, -19573, -14459, -13296, -7813, -3317, 812, 5515, 9568, 13937, 
    18835, 21417, 24573, 26911, 27703, 30342, 30269, 31671, 29897, 28489, 
    28007, 24602, 22466, 19367, 15688, 11686, 8882, 3926, -147, -5006, -9990, 
    -13274, -16932, -20809, -24774, -26767, -28258, -30528, -30465, -31523, 
    -30179, -28936, -27917, -24387, -23544, -20812, -15302, -10982, -8152, 
    -3295, 1464, 3409, 9960, 13298, 16181, 21368, 23140, 25643, 27884, 29632, 
    30383, 31931, 30356, 29205, 29282, 27433, 21977, 19619, 16494, 14318, 
    8350, 3147, 315, -3611, -8150, -12396, -15292, -19706, -22587, -25577, 
    -28248, -29953, -30154, -30547, -30558, -29105, -27179, -27731, -23782, 
    -20249, -15726, -12762, -8852, -4486, 30, 5862, 9051, 12330, 17857, 
    20638, 23655, 24702, 27936, 29008, 30502, 30244, 30027, 29007, 29138, 
    25785, 22485, 19563, 16288, 11837, 9263, 3283, 896, -4374, -8066, -12174, 
    -17159, -20789, -22110, -25537, -26666, -29980, -31551, -30646, -29803, 
    -30338, -28088, -24710, -24123, -19631, -18063, -12352, -9398, -5609, 
    -872, 2502, 7971, 13006, 16094, 21171, 22466, 24865, 27855, 29453, 30909, 
    30656, 30073, 28709, 29307, 26060, 24090, 21134, 16263, 14543, 10868, 
    5291, 751, -4676, -8738, -12313, -16726, -20792, -23299, -26218, -27123, 
    -29532, -30031, -31900, -29329, -30270, -29011, -25803, -25290, -19117, 
    -17146, -12802, -8893, -6837, -1105, 4309, 6757, 12285, 17369, 18196, 
    22599, 25662, 27070, 29705, 30275, 31439, 29375, 30878, 28923, 25854, 
    24354, 21827, 17430, 12620, 9104, 6757, 2719, -2724, -7855, -11416, 
    -14708, -19838, -22629, -24024, -29083, -28143, -29397, -31607, -31769, 
    -30686, -27765, -25968, -23409, -21207, -16280, -12736, -10123, -7426, 
    -995, 3509, 8558, 12777, 15785, 18894, 22883, 26781, 27423, 29874, 30841, 
    30903, 29944, 30334, 28247, 26041, 24195, 21193, 18994, 15921, 8863, 
    6951, 528, -3915, -6576, -11145, -15123, -17600, -23217, -23670, -26092, 
    -29408, -30155, -31375, -30933, -30768, -28858, -26793, -24751, -21566, 
    -18418, -14370, -10478, -5761, -1745, 2906, 5864, 11512, 14514, 17815, 
    22158, 25110, 27910, 28722, 31435, 30727, 30198, 31336, 27997, 26868, 
    25539, 21058, 18177, 13591, 10427, 7519, 491, -2416, -7027, -11174, 
    -14760, -17727, -22118, -24853, -27809, -29374, -29926, -31102, -31417, 
    -30539, -27833, -28045, -24030, -21690, -17815, -14600, -8936, -7654, 
    -2440, 1995, 5107, 11553, 13720, 18453, 22998, 24897, 26692, 28227, 
    29756, 31073, 29412, 31269, 30179, 27391, 24596, 21328, 19296, 14849, 
    11023, 6839, 1904, -2101, -6397, -10448, -14534, -17185, -21421, -24980, 
    -26165, -28708, -30158, -29246, -31759, -28963, -27252, -27474, -25956, 
    -22639, -19403, -14025, -9620, -7932, -3384, 2026, 6105, 9813, 15512, 
    17416, 21339, 24096, 26534, 27960, 29958, 31014, 29735, 29097, 28659, 
    26424, 24073, 21171, 19004, 15411, 11688, 7514, 2225, -1051, -5115, 
    -10870, -13799, -17491, -22348, -24311, -26127, -27922, -29744, -29455, 
    -31411, -30309, -27866, -26920, -26453, -23154, -19750, -14799, -12257, 
    -7487, -2113, 843, 6255, 9633, 12821, 17239, 20889, 23554, 26104, 28676, 
    30355, 30441, 29950, 31394, 28453, 26861, 25490, 21635, 20235, 15897, 
    10074, 7818, 3706, -1802, -3865, -9814, -12970, -16976, -19828, -23816, 
    -26445, -26892, -28843, -30138, -32364, -31568, -29989, -27271, -25452, 
    -22100, -17690, -17049, -10881, -7488, -3546, 859, 6205, 9564, 12819, 
    17373, 19844, 24056, 26396, 29591, 30044, 31465, 30408, 30675, 29519, 
    27852, 24872, 23914, 20355, 14517, 12164, 8217, 3994, -702, -4965, -8684, 
    -12705, -17156, -20884, -23526, -26128, -28828, -29266, -30123, -31540, 
    -31722, -29546, -27774, -24633, -23404, -19576, -15751, -12459, -7975, 
    -3382, 1004, 5306, 9158, 13178, 18246, 20432, 22866, 24960, 29083, 29229, 
    31579, 31651, 29887, 29501, 28155, 25460, 23210, 18290, 16727, 12442, 
    7675, 5688, -1072, -4520, -8326, -11646, -15965, -20754, -23295, -25587, 
    -29112, -29563, -30876, -31157, -31796, -30145, -27780, -25650, -23931, 
    -19778, -15588, -13264, -8867, -3075, -172, 4368, 8425, 12827, 17106, 
    18551, 23412, 25205, 26814, 29053, 29925, 32541, 31431, 29885, 29026, 
    26618, 23528, 21169, 17211, 14369, 9190, 5957, 346, -4488, -8851, -12411, 
    -15098, -20303, -22137, -26311, -28000, -30278, -29501, -30164, -29555, 
    -30349, -28973, -26894, -23259, -20525, -17175, -12634, -9534, -5895, 66, 
    4030, 8773, 12537, 16958, 20116, 23088, 25804, 27338, 30941, 31135, 
    31789, 29589, 29999, 28807, 25845, 22794, 21313, 16357, 13453, 9318, 
    5137, 1209, -3860, -7959, -10592, -16157, -18659, -23838, -25204, -28227, 
    -29990, -29725, -31686, -30243, -28970, -28377, -26574, -24205, -19199, 
    -17311, -13631, -10776, -3706, -870, 4588, 7601, 11075, 15579, 20002, 
    21948, 25123, 27671, 29646, 29250, 30952, 31607, 30240, 28712, 28086, 
    24722, 21332, 18754, 14826, 10500, 5086, 316, -1989, -7564, -11447, 
    -17311, -19942, -23655, -24959, -27274, -27674, -31971, -29586, -30591, 
    -30811, -29333, -26291, -24122, -21376, -17556, -12518, -11470, -7034, 
    -1467, 3421, 7990, 12609, 15445, 19365, 21218, 25194, 27676, 29092, 
    30029, 31108, 31666, 29010, 28430, 27340, 24924, 21815, 17599, 13383, 
    9610, 7085, 1940, -2397, -7264, -10128, -16248, -19093, -22687, -25482, 
    -25691, -27473, -29777, -30495, -30522, -31526, -27694, -27311, -24189, 
    -23258, -17711, -13983, -9590, -5627, -771, 1594, 6499, 12173, 15660, 
    19166, 23234, 23533, 28327, 28622, 30006, 30984, 30983, 28843, 28963, 
    26665, 25670, 22135, 19421, 16219, 9319, 7296, 2182, -3469, -6096, 
    -11303, -13621, -17355, -21364, -25502, -28097, -28423, -29991, -31640, 
    -29804, -30181, -29603, -27338, -23609, -21798, -17547, -13821, -9541, 
    -5305, -1590, 2255, 5750, 9852, 15070, 19022, 21206, 23902, 27536, 28171, 
    30052, 30441, 30258, 30424, 29215, 28531, 24928, 20770, 19762, 14037, 
    9563, 7285, 2039, -3236, -6710, -12305, -15042, -16838, -21189, -24705, 
    -27200, -28264, -30713, -30232, -31001, -30639, -28954, -27476, -25980, 
    -23377, -19067, -15139, -10535, -7000, -4480, 2697, 7098, 10854, 14897, 
    17538, 21511, 25202, 27151, 29058, 29016, 29569, 29362, 29984, 27856, 
    26637, 26270, 20957, 19141, 14265, 12082, 6564, 2504, -2698, -4483, 
    -10105, -14114, -17543, -21152, -24362, -27159, -29684, -30815, -29469, 
    -31264, -29812, -28076, -28026, -24771, -21856, -19474, -15872, -11019, 
    -7638, -2176, -483, 4763, 9549, 15033, 17952, 20820, 25449, 25856, 28500, 
    28531, 31196, 30465, 29829, 28642, 28337, 24970, 22275, 19142, 15374, 
    10939, 6314, 3059, -1864, -6264, -10711, -14835, -16790, -22373, -22655, 
    -26634, -29546, -30236, -31405, -32088, -29741, -27825, -26712, -24246, 
    -23775, -20234, -14316, -11637, -7363, -3713, 1095, 4720, 9956, 13773, 
    17786, 21604, 23304, 27155, 29135, 29568, 31247, 30939, 28934, 29676, 
    27993, 24739, 23391, 19928, 15704, 11631, 8730, 3579, -164, -4922, -9901, 
    -13666, -16923, -21602, -24069, -25620, -28053, -28801, -30335, -30138, 
    -30718, -29818, -29053, -25912, -23484, -21023, -17057, -12836, -9456, 
    -2634, 704, 4254, 8806, 12855, 17407, 19926, 23000, 25473, 28667, 28515, 
    31942, 31332, 30553, 29677, 28428, 24790, 22374, 21169, 17914, 12854, 
    8112, 3787, 722, -4892, -9420, -11226, -15992, -20737, -24009, -25021, 
    -28660, -29434, -29942, -31858, -30724, -29431, -28114, -25165, -23485, 
    -20038, -16300, -12972, -7143, -4007, -340, 4062, 7291, 12317, 16468, 
    19989, 23254, 26755, 28446, 30232, 29229, 31191, 29908, 29873, 26920, 
    25878, 24305, 20543, 17393, 12988, 8667, 4194, 1297, -3517, -8408, 
    -10897, -16438, -21275, -23062, -24740, -26838, -28242, -31823, -31661, 
    -31172, -28710, -27519, -25911, -24151, -20588, -16289, -12739, -9751, 
    -5276, 838, 4318, 8701, 12640, 15688, 19016, 23165, 25845, 27948, 29557, 
    30847, 30231, 30538, 31543, 27893, 26108, 23137, 19514, 15458, 14201, 
    8807, 4599, 456, -2028, -6957, -12054, -16744, -19262, -22301, -26161, 
    -26505, -30343, -30305, -31404, -31506, -30360, -28004, -26516, -23644, 
    -20696, -17414, -14227, -11055, -4805, -2178, 4136, 7809, 10572, 16181, 
    18872, 21805, 26094, 28499, 29235, 29191, 30961, 31013, 31084, 27947, 
    26009, 23871, 20864, 18459, 14383, 10197, 4024, 886, -3394, -6292, 
    -11575, -15252, -20162, -22976, -25390, -25868, -29276, -31071, -31208, 
    -30084, -28313, -30026, -25692, -24162, -22615, -16405, -14659, -10581, 
    -7038, -1463, 2515, 6992, 10012, 16401, 19694, 21214, 25487, 28738, 
    28203, 30052, 31112, 30604, 30203, 27592, 25316, 25392, 19893, 16959, 
    14143, 10804, 6031, 2348, -2907, -7469, -11657, -16406, -19208, -22774, 
    -26420, -27058, -29629, -31415, -30463, -29443, -29866, -29062, -26905, 
    -25061, -21472, -18632, -14214, -10124, -6741, -2115, 2644, 6579, 11037, 
    16322, 18894, 23073, 25573, 27359, 28839, 30343, 31112, 30561, 30015, 
    28889, 27064, 24175, 22364, 18845, 13599, 11031, 6034, 2248, -2551, 
    -6690, -10631, -14149, -17261, -20385, -25626, -26829, -29352, -30115, 
    -31289, -30410, -31692, -28892, -27737, -24226, -21567, -17856, -14604, 
    -10767, -6784, -1537, 2147, 6384, 10090, 15341, 17400, 21008, 24389, 
    27319, 28174, 30322, 31385, 31048, 30517, 28725, 25631, 23364, 21123, 
    17840, 14532, 9673, 5351, 1522, -604, -6641, -9810, -14687, -17676, 
    -22446, -23960, -27168, -27824, -30041, -30802, -30547, -29351, -30117, 
    -27222, -25788, -22103, -19262, -14275, -12303, -5320, -2246, 2281, 6765, 
    9426, 13576, 17693, 21552, 24412, 25963, 29990, 29785, 31074, 31442, 
    31528, 29097, 27351, 25797, 22780, 19792, 14258, 11029, 7264, 2311, 
    -1154, -5001, -11110, -13094, -17864, -21860, -24085, -26953, -28566, 
    -29567, -31363, -30897, -31191, -30800, -27823, -24966, -22811, -18209, 
    -15727, -11231, -6752, -1814, 1066, 5288, 10491, 14587, 17429, 21872, 
    22567, 26016, 29223, 29593, 30197, 30184, 31169, 29409, 27865, 24605, 
    23378, 19932, 16518, 12114, 8720, 3152, -2739, -4811, -9311, -15093, 
    -16852, -21282, -24095, -25780, -28841, -30033, -31871, -31517, -29959, 
    -29552, -28209, -24525, -22299, -20355, -15851, -10880, -5991, -4713, 
    1521, 4578, 8776, 14065, 18147, 22008, 23058, 26679, 28923, 30778, 31277, 
    31888, 29711, 28009, 27878, 24428, 22423, 18489, 16614, 12683, 7083, 
    3440, -1047, -5892, -10088, -12698, -17525, -20161, -25341, -26300, 
    -29177, -30080, -31225, -31420, -31283, -29104, -28142, -26434, -22709, 
    -19445, -16176, -12575, -8187, -3534, 1886, 4142, 9574, 13254, 17934, 
    21036, 22492, 25895, 29530, 29281, 30829, 30662, 30986, 31008, 28967, 
    27151, 22850, 18342, 17147, 13132, 8356, 3501, -1851, -4538, -9647, 
    -12793, -15739, -21718, -23244, -25410, -27818, -30183, -30297, -30912, 
    -30140, -28703, -28044, -25960, -23209, -20330, -16107, -13148, -8109, 
    -5377, -1013, 5295, 8247, 12462, 15263, 18617, 21747, 25999, 27357, 
    29621, 31678, 29858, 29711, 29516, 26998, 24947, 22716, 20232, 16078, 
    11894, 9626, 4186, 568, -3386, -7892, -11793, -17120, -19020, -23854, 
    -25337, -29287, -29916, -30530, -30556, -30587, -30573, -27097, -25687, 
    -23672, -19693, -18328, -12633, -8910, -4341, -1133, 3959, 6944, 11884, 
    16243, 19932, 23734, 25312, 28156, 28944, 29557, 30240, 29426, 30832, 
    28337, 25845, 23892, 21384, 15664, 14013, 8276, 5964, -177, -4299, -8464, 
    -11609, -15498, -18461, -23992, -25811, -28138, -29561, -31064, -30609, 
    -30989, -29426, -27665, -26683, -23037, -20312, -17169, -12720, -10266, 
    -4997, -252, 4322, 7514, 11899, 16098, 18748, 22917, 24752, 27157, 29737, 
    30318, 31283, 30765, 30796, 28678, 26370, 22795, 21410, 17318, 13988, 
    10663, 5617, 1896, -3681, -7622, -12767, -16522, -19048, -20992, -24447, 
    -28200, -30289, -30244, -30934, -31101, -29609, -28535, -26010, -23957, 
    -20525, -18586, -13780, -8662, -5559, -241, 2911, 7812, 10978, 15170, 
    18869, 23466, 24287, 27468, 28714, 29713, 30029, 29010, 30413, 30252, 
    26422, 23948, 21901, 17908, 13085, 9249, 6009, 565, -1868, -8853, -11894, 
    -15094, -17420, -21019, -25440, -27323, -28973, -31485, -31427, -29937, 
    -29734, -28361, -28299, -24346, -21706, -17855, -14293, -11772, -6797, 
    -1661, 1274, 7246, 10854, 14973, 18193, 21986, 26641, 28877, 28565, 
    29634, 31125, 30538, 30563, 29376, 26212, 23890, 21650, 17252, 14792, 
    9755, 5974, 2865, -3300, -6891, -9425, -16078, -19193, -22592, -25381, 
    -27861, -29049, -30217, -29017, -29938, -31103, -27657, -26726, -24956, 
    -22579, -18557, -14663, -10564, -5878, -886, 2665, 5996, 9545, 15727, 
    17510, 20820, 24989, 27785, 27826, 30528, 31109, 29967, 30145, 28816, 
    26563, 25719, 23031, 17342, 13981, 11208, 7192, 1586, -1626, -7195, 
    -10011, -14670, -17745, -21973, -24854, -26279, -28535, -30430, -30705, 
    -31923, -31076, -29329, -27232, -23838, -21829, -17087, -13740, -10207, 
    -6263, -3274, 465, 5705, 11410, 13401, 17203, 21445, 25133, 28353, 27755, 
    31114, 29413, 29519, 29555, 30190, 28757, 23974, 22368, 19133, 16645, 
    10738, 6975, 3664, -2209, -5109, -11761, -14167, -18199, -22928, -24955, 
    -26552, -27973, -28698, -30179, -30509, -30517, -29967, -26580, -24883, 
    -21181, -18725, -15545, -10910, -6692, -3769, 1078, 5780, 9468, 13736, 
    17297, 21268, 24447, 25926, 27063, 29553, 31122, 30734, 29783, 29812, 
    28042, 25971, 23129, 18872, 16417, 11805, 8060, 3639, -450, -6298, -9546, 
    -15083, -17168, -21720, -24292, -24917, -29133, -29773, -31527, -29472, 
    -30081, -29132, -27833, -25486, -23136, -19227, -17049, -10660, -8158, 
    -2983, 1676, 5061, 10031, 12794, 17081, 21610, 23370, 26913, 27826, 
    29955, 31727, 31496, 31036, 29563, 28045, 26017, 23362, 19442, 17237, 
    12486, 8479, 5241, -1374, -4943, -8556, -14480, -16061, -19776, -24270, 
    -26177, -28390, -29621, -30718, -30369, -30869, -29401, -27152, -26055, 
    -23364, -19921, -17818, -12291, -7746, -4335, 464, 4915, 10166, 11956, 
    16121, 19620, 24753, 25419, 29235, 28980, 30582, 32316, 30862, 27872, 
    27490, 25747, 22096, 19899, 16666, 12721, 8454, 3606, 1086, -5167, -9132, 
    -13524, -17344, -21307, -23171, -27493, -28048, -30043, -30573, -31366, 
    -31674, -29115, -26359, -26429, -23019, -19991, -16524, -13582, -8534, 
    -3878, 650, 4108, 7751, 13015, 16787, 21129, 23003, 26029, 26708, 29146, 
    30240, 30446, 29591, 29614, 27796, 26817, 23298, 20019, 15918, 13294, 
    7037, 3941, -358, -4061, -9635, -11953, -15487, -19751, -24345, -25942, 
    -26805, -30463, -30981, -30450, -30608, -29234, -28483, -24697, -24046, 
    -20887, -15747, -11437, -8568, -3965, -1631, 4818, 9070, 12805, 16559, 
    19938, 23834, 25314, 27997, 28345, 29484, 31011, 31357, 28341, 28550, 
    26956, 23802, 20516, 15816, 12384, 10001, 4712, 1166, -4373, -7805, 
    -12740, -15591, -19687, -23502, -24645, -28178, -29914, -31251, -31057, 
    -31102, -29008, -27969, -26227, -24980, -19568, -17505, -14303, -9792, 
    -4051, -721, 2632, 8730, 12850, 17311, 19401, 22725, 23913, 28003, 28297, 
    29479, 30444, 31074, 28831, 28293, 25271, 22135, 20791, 18074, 13298, 
    9961, 5619, 1260, -2408, -6528, -11694, -15576, -20346, -21745, -25760, 
    -28027, -29523, -30993, -30696, -30893, -29914, -28582, -25995, -24989, 
    -19731, -17362, -14295, -9941, -5598, -307, 3280, 6009, 11074, 14722, 
    18532, 21761, 24564, 27788, 28917, 31668, 32482, 31999, 30271, 28747, 
    27047, 24909, 20112, 18328, 14221, 8825, 5353, 1096, -3612, -6465, 
    -12796, -16071, -19072, -21620, -23980, -27850, -29624, -29584, -31450, 
    -30937, -30349, -28750, -26350, -24540, -20188, -18441, -14199, -10491, 
    -5814, -1683, 3852, 7128, 10501, 16318, 19002, 22654, 25726, 27864, 
    28020, 29327, 30613, 29763, 30347, 28805, 26722, 23570, 22184, 20065, 
    14969, 10560, 6666, 2392, -1735, -5008, -11016, -15226, -19140, -23636, 
    -23820, -27178, -29334, -29958, -29563, -29270, -30540, -28780, -26130, 
    -24588, -23171, -16761, -14154, -9532, -7407, -2224, 2736, 7576, 9960, 
    14335, 18050, 21242, 24457, 28744, 30277, 29763, 30881, 30931, 28844, 
    29708, 27247, 25088, 23686, 18901, 15488, 11574, 5392, 3840, -3166, 
    -5437, -10563, -15693, -18615, -23263, -24351, -26161, -28530, -29304, 
    -30807, -30878, -30157, -28837, -27762, -24309, -21749, -20130, -16324, 
    -10684, -7455, -4055, 1276, 5081, 9899, 14475, 16458, 20921, 24626, 
    25198, 30398, 31315, 31430, 30218, 30754, 30024, 27920, 25790, 23688, 
    19426, 15813, 11948, 8122, 2883, -1219, -5181, -8666, -14582, -17218, 
    -22042, -25822, -26712, -28393, -29676, -31319, -30865, -30306, -29353, 
    -27331, -25165, -22708, -18891, -16428, -13057, -6206, -3763, 1030, 4285, 
    9886, 15560, 18252, 20330, 23263, 27210, 26936, 30942, 30714, 30020, 
    31418, 29854, 27235, 25538, 22894, 20459, 15530, 12600, 6668, 2845, 
    -1465, -3998, -8971, -13348, -17810, -21680, -25069, -26366, -28523, 
    -29666, -30046, -31142, -30166, -28036, -26543, -23773, -23276, -19400, 
    -15210, -11428, -8574, -3990, 594, 5418, 9543, 12047, 18280, 21937, 
    23632, 26048, 27827, 31361, 29394, 32222, 30319, 28718, 27217, 25851, 
    22375, 19246, 16649, 11969, 8371, 2061, -862, -4878, -10177, -12618, 
    -18681, -20563, -23109, -26203, -28459, -30156, -30004, -30387, -29959, 
    -30975, -27666, -26653, -23313, -19627, -16787, -12430, -8634, -4132, 
    1611, 4114, 8989, 13540, 18432, 20686, 22556, 25924, 28242, 28239, 31759, 
    31466, 30797, 30733, 27550, 25607, 23757, 21025, 16268, 11917, 9582, 
    5864, -449, -5707, -8740, -13315, -17952, -20493, -23474, -25691, -27704, 
    -28885, -30304, -30043, -30505, -29231, -27017, -26586, -24383, -20282, 
    -17752, -12369, -7655, -5099, -1226, 4372, 8793, 13272, 16181, 19387, 
    24454, 24630, 28757, 29952, 29157, 31274, 29563, 29869, 28934, 25991, 
    25062, 20871, 16246, 13420, 7519, 3094, 931, -5015, -7928, -12470, 
    -16550, -20288, -23275, -25750, -28224, -29142, -30326, -31087, -31321, 
    -28411, -28355, -26103, -23489, -20832, -16223, -12471, -9273, -4890, 
    -1519, 3818, 9439, 10548, 15961, 18345, 21867, 24794, 27776, 28259, 
    31522, 32449, 30980, 29719, 28166, 27152, 23807, 20050, 16842, 13752, 
    9700, 4323, 762, -4331, -7891, -13097, -15815, -19595, -22234, -24560, 
    -27674, -29461, -30505, -31278, -29217, -28173, -27646, -26477, -24777, 
    -21867, -17464, -13186, -9351, -4337, 84, 3726, 8373, 11293, 14776, 
    20042, 22137, 27150, 27080, 28755, 30416, 30729, 31712, 29693, 28311, 
    26355, 23525, 20510, 17646, 14800, 9832, 5722, 81, -3253, -7895, -11245, 
    -15606, -19303, -22478, -25490, -26731, -29396, -31626, -30670, -30968, 
    -29455, -27423, -26923, -24517, -20158, -18628, -14882, -9609, -5567, 
    -1957, 3036, 8205, 10641, 16497, 17804, 21114, 23324, 27159, 28343, 
    31530, 29497, 30160, 30228, 28940, 25317, 24247, 22768, 18008, 15380, 
    9897, 4929, 2471, -2772, -7099, -10733, -16777, -18548, -21073, -24158, 
    -27213, -27977, -30765, -31780, -31492, -30495, -28336, -28154, -23784, 
    -21705, -17311, -15056, -10400, -5139, -894, 1579, 6964, 11969, 14566, 
    18960, 23049, 25075, 27896, 27213, 30343, 30621, 29563, 29691, 27532, 
    27403, 24144, 23319, 18942, 14700, 10605, 6721, 2845, -3253, -5815, 
    -11185, -16359, -18045, -22438, -25111, -26761, -30439, -29334, -32464, 
    -31400, -31138, -28952, -26729, -24127, -22219, -18632, -15819, -11713, 
    -7068, -1765, 2823, 7263, 12376, 15029, 18910, 23035, 24995, 26819, 
    28695, 30059, 30646, 30924, 28587, 28184, 26495, 26545, 21264, 18711, 
    13419, 11130, 6807, 988, -2893, -7255, -10123, -14900, -18052, -20185, 
    -24013, -27639, -30167, -29969, -30945, -29739, -31784, -29935, -27364, 
    -23734, -23088, -19504, -14332, -10796, -7215, -3241, 2549, 5580, 11038, 
    14380, 19435, 20097, 24780, 26598, 28864, 29896, 32046, 29301, 31338, 
    28440, 26528, 25056, 20574, 17632, 14212, 12202, 6237, 2990, -2513, 
    -6155, -9468, -14556, -16862, -20237, -23365, -26575, -28062, -30030, 
    -31332, -30850, -30883, -28984, -28520, -25735, -22552, -18619, -15117, 
    -9977, -7294, -3236, 2258, 6295, 9283, 13857, 19285, 20056, 24129, 26480, 
    29015, 28446, 30656, 31026, 30079, 30908, 27454, 25147, 22156, 18531, 
    15999, 10975, 7837, 2726, -1113, -5099, -8890, -13810, -17503, -19737, 
    -23440, -26472, -29047, -31104, -30161, -30315, -30697, -29869, -27914, 
    -25610, -22914, -19188, -15663, -13306, -8003, -3099, 776, 4160, 10161, 
    13797, 17914, 22368, 22760, 26872, 28213, 30420, 29859, 29598, 30729, 
    29131, 28249, 24424, 23188, 20843, 15493, 12876, 6320, 3672, -1612, 
    -6066, -9389, -12359, -17481, -19490, -23423, -27209, -27443, -31531, 
    -30677, -30559, -29923, -28636, -28526, -24359, -22691, -20462, -15810, 
    -12019, -8446, -2558, 862, 5134, 9802, 11419, 16755, 20067, 21943, 25646, 
    27007, 29622, 30924, 31640, 31929, 29880, 27466, 25454, 23766, 20106, 
    16020, 13835, 7074, 3316, 390, -4396, -9559, -12626, -16462, -21332, 
    -23021, -24735, -27759, -29116, -30357, -31655, -30431, -29432, -27580, 
    -26599, -22855, -19502, -17913, -13258, -8018, -4850, -164, 4003, 7671, 
    11691, 16148, 20627, 23609, 25622, 26777, 30249, 30667, 31826, 30714, 
    30281, 27207, 24801, 23330, 20533, 16411, 13097, 9468, 4287, 171, -2685, 
    -8201, -12030, -14743, -20154, -24596, -24212, -27130, -28225, -30301, 
    -30412, -28918, -29738, -27395, -27498, -23839, -19213, -15861, -14855, 
    -8743, -4889, -904, 4243, 6664, 12489, 15665, 19673, 23136, 26027, 28598, 
    30838, 30261, 32028, 29624, 29428, 28814, 26816, 22438, 21851, 16916, 
    11986, 9122, 3627, 10, -3785, -7396, -13231, -16099, -19747, -24088, 
    -26470, -27405, -29864, -29588, -29630, -30451, -29400, -29261, -27387, 
    -23039, -21377, -17553, -13619, -10357, -5077, -388, 4372, 8791, 12545, 
    15862, 20851, 21079, 25116, 27733, 29069, 29978, 30820, 29739, 29792, 
    28092, 27804, 24062, 21200, 16854, 14080, 11339, 4876, 1465, -2348, 
    -6356, -11554, -15548, -19967, -21870, -24645, -28247, -28085, -31740, 
    -32338, -31364, -30443, -29693, -27448, -22501, -20103, -17407, -12206, 
    -9730, -6378, -1174, 3256, 8470, 11176, 15710, 20240, 22771, 26199, 
    27054, 29978, 29261, 30004, 31004, 30381, 29478, 26907, 24674, 20374, 
    17590, 15222, 9073, 6383, 1095, -4063, -7428, -12025, -14835, -19940, 
    -22433, -24635, -26586, -30195, -30323, -30645, -29895, -29568, -28872, 
    -27796, -23513, -21103, -17888, -14777, -10513, -5685, -1253, 2967, 6680, 
    11389, 15329, 17492, 21873, 23756, 28633, 30361, 30194, 30906, 32043, 
    31055, 28623, 26799, 24280, 22864, 17283, 14396, 10950, 6588, 3157, 
    -2627, -7018, -11936, -15056, -19809, -22894, -23278, -28197, -28858, 
    -30006, -32043, -31438, -28650, -29829, -26082, -23601, -22511, -18496, 
    -13439, -9947, -7278, -1989, 1460, 7151, 10846, 14361, 18671, 20372, 
    25977, 26764, 29918, 30788, 30215, 29533, 30553, 29476, 28035, 24313, 
    22633, 18727, 14410, 10486, 6913, 2686, -1887, -6457, -9144, -13680, 
    -19075, -21417, -25894, -26733, -29117, -29237, -31735, -30981, -30180, 
    -28422, -26280, -25698, -23451, -18863, -16000, -11418, -5638, -2945, 
    2248, 6242, 11781, 15702, 17298, 22823, 24349, 27721, 28274, 31364, 
    30854, 30647, 29830, 29774, 26840, 25030, 21564, 19217, 14332, 11177, 
    6349, 3059, -1558, -5852, -8929, -15632, -17376, -22243, -25431, -25997, 
    -29238, -28658, -32138, -31011, -29276, -29043, -26582, -26392, -23354, 
    -18422, -15874, -12229, -7577, -3010, 2188, 5644, 9052, 13177, 17593, 
    20395, 23011, 26263, 27374, 28804, 29071, 30065, 29117, 29388, 27922, 
    26325, 23101, 19392, 15014, 12257, 9197, 3918, -920, -4245, -9931, 
    -13798, -17688, -21766, -24865, -25787, -27317, -30326, -29790, -30736, 
    -29526, -27778, -27222, -26070, -23697, -20466, -14965, -11307, -6312, 
    -3982, 206, 5174, 8798, 13728, 18416, 19136, 22914, 26362, 27547, 29738, 
    32123, 31170, 30285, 28457, 27666, 24158, 23448, 19882, 16392, 13386, 
    7048, 4175, -1040, -4156, -10048, -14692, -16414, -20356, -23157, -25687, 
    -28382, -29591, -31932, -29433, -30162, -29102, -29068, -25915, -22458, 
    -21136, -15952, -13495, -8458, -4899, -330, 4789, 9692, 12469, 16131, 
    21080, 22991, 26466, 28919, 30228, 30780, 31814, 30980, 28911, 27946, 
    25930, 23682, 21410, 18153, 13016, 6912, 4497, 283, -4955, -8891, -14090, 
    -15329, -19136, -23067, -25496, -26678, -28886, -30788, -32178, -31208, 
    -30006, -28797, -25400, -22678, -20283, -16969, -12949, -7117, -4629, 
    569, 4175, 7015, 11944, 16706, 20448, 22785, 25637, 26504, 29910, 29639, 
    30932, 29925, 29696, 28058, 26518, 23867, 20475, 17997, 12117, 8331, 
    3511, -523, -4478, -8817, -12007, -16521, -19169, -23914, -26115, -27367, 
    -30604, -30828, -30839, -29382, -27930, -28178, -26112, -23989, -19206, 
    -18478, -13976, -9860, -4963, -1019, 3806, 7933, 13719, 16236, 18790, 
    24588, 25340, 28144, 30153, 30334, 30815, 29776, 31224, 27822, 26565, 
    24474, 20130, 17183, 13526, 11127, 5170, 1013, -3080, -8647, -12637, 
    -15889, -21136, -22598, -25100, -25899, -30453, -29870, -32170, -30064, 
    -29209, -28294, -26313, -24369, -20810, -16969, -13440, -8891, -6398, 
    -333, 3543, 7383, 11392, 15950, 20193, 21488, 24894, 27255, 29748, 29768, 
    31107, 29803, 29608, 28280, 26972, 25363, 20822, 17804, 13037, 9011, 
    6183, 1549, -2354, -7603, -13088, -16537, -19684, -22867, -24352, -28712, 
    -28809, -29796, -30048, -30567, -28826, -28118, -25744, -24314, -20547, 
    -16692, -12858, -10004, -4429, -988, 2729, 8205, 12303, 15378, 18241, 
    21871, 26160, 27547, 29841, 31501, 30097, 31669, 29872, 29948, 26775, 
    24271, 22404, 17643, 13313, 9975, 6300, 830, -2373, -5844, -10115, 
    -15468, -19612, -23715, -24714, -27780, -28935, -28354, -30650, -31116, 
    -29507, -29428, -26983, -23732, -21168, -18517, -15384, -9544, -5738, 
    -1407, 3654, 5780, 10158, 16667, 17476, 22887, 24160, 26474, 30615, 
    29421, 29418, 31119, 29494, 30569, 26405, 24553, 21796, 18141, 14009, 
    11444, 6450, 2367, -1380, -7417, -11219, -16016, -19538, -21844, -24909, 
    -26157, -27915, -28917, -29561, -30767, -30268, -28580, -27616, -25134, 
    -22666, -18999, -13608, -12675, -7965, -1193, 2892, 5241, 9633, 14821, 
    17428, 22305, 24386, 27322, 29412, 29807, 30470, 30579, 28687, 28246, 
    26520, 24924, 21801, 18286, 15008, 11904, 6379, 1978, -1777, -6219, 
    -11244, -13548, -17385, -22404, -24869, -27093, -29455, -29356, -30140, 
    -31584, -30915, -28230, -28412, -23726, -20521, -17733, -14735, -11324, 
    -7154, -2140, 1572, 7089, 11638, 14665, 19506, 22121, 24657, 27526, 
    30060, 30152, 30365, 29868, 28544, 29884, 28348, 26216, 21937, 19656, 
    15281, 10361, 5706, 3041, -1061, -5476, -10288, -14723, -18351, -21065, 
    -23716, -27516, -29966, -30816, -31318, -29685, -29321, -30083, -28381, 
    -25197, -21888, -19322, -15726, -11186, -7643, -1962, 1576, 5938, 9749, 
    14272, 17830, 21947, 25643, 27824, 28348, 30526, 29062, 30045, 28670, 
    30022, 27671, 24050, 22422, 19346, 15142, 13107, 6417, 4061, -748, -4673, 
    -8756, -14435, -18046, -21548, -24062, -27567, -28433, -29525, -31387, 
    -30122, -30814, -28127, -28115, -25097, -23418, -20316, -15870, -10638, 
    -7170, -2116, 1240, 4313, 9471, 13182, 16812, 21643, 23421, 27376, 28155, 
    28921, 30148, 30934, 32122, 29964, 27787, 24338, 21802, 19862, 16095, 
    10833, 9066, 3245, -208, -6390, -8758, -12160, -15301, -20610, -25124, 
    -25033, -29030, -28487, -30370, -31126, -30857, -29594, -27759, -25664, 
    -24542, -19943, -16202, -11223, -7723, -2506, 2228, 4589, 8157, 12365, 
    17127, 21505, 22890, 26140, 29854, 29713, 29520, 30107, 30420, 29247, 
    26708, 25247, 21895, 19134, 16277, 11629, 8474, 4515, -730, -4221, -8179, 
    -13194, -17684, -20727, -22167, -25865, -26695, -28292, -30914, -30225, 
    -29302, -29724, -29364, -25896, -23752, -19668, -15553, -13091, -7454, 
    -4427, 379, 4328, 9407, 11721, 16767, 21989, 21592, 26768, 27964, 30241, 
    30751, 31093, 30841, 30192, 29143, 25925, 22520, 21394, 17110, 13228, 
    8374, 3638, 1597, -4178, -8891, -12916, -16396, -21871, -21976, -25987, 
    -28200, -30092, -29946, -30858, -31527, -29783, -28065, -25733, -23142, 
    -21300, -16794, -12854, -10556, -4322, -614, 2798, 7853, 12983, 15500, 
    19032, 24105, 24362, 27743, 30250, 30839, 31680, 30732, 30353, 28830, 
    26912, 25459, 20364, 17776, 13669, 8380, 4926, 1164, -3853, -7906, 
    -10685, -16076, -19622, -23830, -24706, -28993, -29309, -30270, -30020, 
    -30637, -30319, -29019, -24884, -25661, -19742, -17997, -13583, -8490, 
    -5458, -1273, 3102, 6465, 12349, 16872, 20306, 22939, 24889, 28263, 
    29170, 30725, 31146, 30224, 29977, 29270, 26230, 24330, 20842, 17005, 
    13673, 9883, 6378, 614, -3154, -6553, -12558, -14568, -19294, -22341, 
    -25003, -27449, -29310, -29304, -31676, -30938, -28782, -29826, -26034, 
    -23122, -19559, -17724, -13941, -10272, -4875, -1404, 2187, 6203, 12132, 
    14203, 18188, 21683, 26188, 26366, 30679, 29789, 29257, 30857, 29301, 
    28985, 26611, 25076, 20909, 18242, 14647, 11769, 5698, 994, -3862, -6494, 
    -11158, -14254, -19469, -22440, -24594, -27967, -28313, -29701, -29550, 
    -29160, -29264, -28722, -26870, -25544, -20939, -18823, -13308, -9110, 
    -6059, -1469, 1721, 6804, 12425, 14951, 18632, 22693, 23747, 27915, 
    27356, 29559, 30580, 31748, 29234, 27655, 26718, 23188, 20885, 18795, 
    16223, 11439, 5853, 1074, -3849, -6270, -10764, -14450, -19326, -21813, 
    -24948, -27030, -30131, -29072, -31239, -31158, -29451, -29357, -26202, 
    -24850, -21673, -19129, -13542, -9786, -6834, -2519, 2947, 5162, 12043, 
    14071, 17072, 22070, 23794, 25530, 29552, 29176, 30844, 31155, 29600, 
    27917, 27401, 25183, 22063, 17934, 15223, 11236, 6516, 2058, -1492, 
    -6060, -10086, -14011, -18688, -21023, -23335, -26992, -28182, -29619, 
    -32240, -30185, -29401, -28575, -26682, -25184, -21577, -18190, -15375, 
    -9873, -7188, -2722, 1057, 4882, 10903, 13525, 18540, 21633, 22821, 
    28290, 27679, 30096, 30002, 29440, 30813, 28853, 25840, 24846, 23017, 
    18654, 15839, 10715, 6690, 2066, -579, -7141, -10835, -14396, -18557, 
    -22466, -24771, -26993, -28861, -28831, -31323, -32356, -31102, -27995, 
    -26337, -25084, -23512, -18637, -17246, -10590, -5914, -4072, 2378, 5908, 
    9982, 14089, 16479, 20983, 23592, 26834, 29823, 30557, 31227, 29649, 
    31140, 28763, 26656, 25681, 21262, 19263, 14016, 12091, 8798, 3736, 
    -2096, -4020, -11185, -15478, -18228, -20088, -23341, -26073, -28737, 
    -30101, -30802, -32011, -28812, -30536, -28106, -25432, -23226, -20297, 
    -14614, -12597, -7467, -4068, 2243, 5326, 10778, 12527, 17734, 20741, 
    23432, 25988, 28909, 29316, 29677, 31743, 31281, 29357, 27297, 25908, 
    22194, 20005, 16377, 11545, 8675, 3863, -387, -6235, -7544, -11819, 
    -16824, -18751, -22918, -26700, -27252, -30499, -29549, -30363, -30960, 
    -27713, -26511, -24269, -22999, -20587, -17260, -12276, -9845, -3412, 
    1200, 5456, 8465, 11865, 16498, 19452, 23400, 26376, 29613, 28882, 29951, 
    30263, 30674, 29763, 28199, 26316, 24220, 21445, 15865, 13414, 8394, 
    3908, 772, -4266, -8429, -12757, -17193, -19090, -23343, -27198, -28198, 
    -30416, -32017, -29333, -30062, -30166, -27874, -25715, -22461, -21248, 
    -16523, -14038, -8536, -4464, -602, 5917, 7891, 11738, 16375, 19750, 
    23405, 24980, 28150, 28538, 31954, 30908, 31103, 29756, 26911, 25974, 
    22862, 20404, 17461, 12752, 9184, 4505, 754, -3948, -8036, -12442, 
    -16746, -20350, -22667, -26270, -28126, -28142, -30560, -29791, -29501, 
    -30655, -28242, -26043, -23493, -20008, -17185, -12040, -8708, -4375, 
    -1781, 4913, 7967, 11890, 15047, 18464, 22628, 24942, 28514, 30490, 
    29866, 31673, 30082, 30575, 29212, 25214, 24046, 20983, 18702, 12427, 
    7736, 5276, 589, -3079, -6938, -12855, -16239, -19830, -23755, -26082, 
    -28525, -28537, -29038, -32193, -31911, -29739, -28755, -25502, -23965, 
    -22165, -17343, -13171, -10672, -6179, -473, 1976, 8923, 11258, 17564, 
    19570, 23378, 25427, 29071, 28059, 30095, 30691, 31261, 29390, 28673, 
    26196, 23910, 19800, 16917, 14447, 9511, 4191, 957, -3493, -8005, -12298, 
    -15449, -20579, -23878, -26112, -29064, -28861, -29986, -29954, -29980, 
    -28910, -28151, -27037, -23596, -21564, -17930, -13917, -9451, -7061, 
    -1435, 2188, 7400, 10484, 14209, 19452, 20833, 24623, 28093, 30264, 
    29834, 29717, 29078, 30818, 28468, 27146, 25038, 21873, 17938, 12749, 
    10492, 6134, -272, -4181, -6963, -11890, -15155, -18196, -22298, -25271, 
    -27160, -28424, -30053, -30506, -30800, -30000, -29374, -25758, -24506, 
    -22870, -19123, -14601, -10366, -6542, -2241, 2385, 6610, 10055, 16156, 
    18882, 21463, 24182, 26875, 29608, 30144, 31282, 29841, 28769, 29665, 
    27795, 23035, 21011, 19032, 14647, 11453, 5745, 651, -2668, -6778, 
    -10866, -13797, -19230, -20554, -24482, -25793, -28984, -29512, -32140, 
    -30158, -31253, -29166, -28054, -24439, -21572, -19166, -14698, -10134, 
    -7363, -3283, 2193, 6559, 11821, 14864, 18959, 20148, 23467, 28478, 
    29601, 29105, 31488, 29586, 30563, 28768, 26518, 23753, 22488, 18596, 
    13221, 12339, 6677, 2148, -2714, -5317, -10146, -14312, -19223, -21288, 
    -23952, -28209, -27879, -28661, -30496, -30070, -29656, -27600, -26509, 
    -24110, -21398, -17575, -14463, -11495, -5222, -2732, 928, 5486, 10342, 
    12870, 16577, 21505, 24977, 26256, 29040, 30026, 29798, 30295, 30065, 
    28338, 26743, 25001, 22457, 19491, 15573, 11972, 7345, 1140, -1123, 
    -6809, -10572, -13977, -18198, -21737, -24779, -25323, -29125, -28607, 
    -31358, -31542, -31559, -28357, -27745, -25303, -21124, -20777, -15094, 
    -11100, -6183, -3601, 1800, 4646, 8985, 13306, 18829, 19932, 23728, 
    26905, 27193, 29746, 30567, 30394, 28869, 29668, 27297, 25024, 23834, 
    20264, 16174, 13105, 7552, 4191, -293, -4636, -9650, -14179, -17171, 
    -19365, -25241, -26396, -29726, -30574, -30901, -29755, -30735, -27841, 
    -28310, -25571, -23241, -19074, -15496, -11233, -7647, -3854, 2039, 4889, 
    8344, 14754, 16121, 19960, 23370, 26347, 28489, 29754, 30487, 32215, 
    31777, 28861, 27836, 26575, 22511, 19467, 16383, 11452, 6879, 3152, 112, 
    -5431, -10486, -13165, -17111, -19925, -23393, -26012, -27873, -29880, 
    -29463, -31117, -31626, -28111, -26012, -25085, -23667, -20449, -15370, 
    -12549, -7024, -4463, 11, 4653, 9718, 13382, 16986, 21149, 24592, 25980, 
    29227, 29352, 30812, 31527, 32045, 27945, 27940, 26908, 22263, 21451, 
    16248, 13370, 8393, 2825, -636, -5087, -9788, -12897, -18370, -18799, 
    -24028, -26019, -29657, -29828, -30252, -29990, -30321, -28897, -27868, 
    -26195, -23349, -20742, -16826, -13166, -8950, -4339, -85, 5274, 8383, 
    12369, 18272, 19987, 22779, 27030, 27135, 28028, 29661, 31811, 31143, 
    29974, 29633, 26733, 23884, 20279, 17520, 14193, 8279, 3417, -876, -4087, 
    -9710, -10826, -16727, -19746, -22821, -26803, -29080, -28874, -30772, 
    -30589, -30991, -29831, -27416, -25699, -24775, -20939, -16799, -14047, 
    -9652, -5498, -1519, 4133, 7757, 13369, 15681, 21017, 22653, 26386, 
    28483, 29304, 29373, 30853, 30812, 29753, 27723, 25054, 23563, 22033, 
    16422, 13007, 8312, 3903, 634, -3914, -6828, -11614, -15454, -21105, 
    -22040, -24922, -27413, -29666, -32220, -30524, -31736, -29292, -29207, 
    -27034, -23156, -19682, -17384, -13210, -9036, -5078, -1575, 4812, 7820, 
    11353, 15730, 20276, 23298, 25536, 27522, 30491, 31733, 30176, 30468, 
    29336, 28840, 27153, 24385, 19990, 17335, 15278, 10334, 4894, -573, 
    -3944, -8844, -12110, -16502, -19970, -21478, -24797, -27769, -29122, 
    -29927, -30060, -30323, -29542, -29019, -25751, -25297, -19882, -17291, 
    -14050, -9622, -5342, -1924, 3452, 8582, 10358, 16164, 17388, 22118, 
    25425, 28161, 29436, 30761, 30382, 29951, 29728, 27217, 26795, 24011, 
    21781, 16846, 13614, 10270, 7119, 947, -2700, -7041, -10131, -16043, 
    -18787, -21536, -25653, -28234, -30389, -29577, -30231, -30438, -30699, 
    -29596, -26562, -24256, -20257, -19284, -14669, -10164, -6693, -1997, 
    1815, 7257, 11540, 15008, 19415, 22197, 24707, 26329, 28848, 30269, 
    29882, 31776, 29859, 28564, 26855, 23255, 21658, 18388, 14679, 9122, 
    5575, 728, -1543, -5612, -11817, -16057, -16914, -20968, -24474, -27134, 
    -28062, -30837, -29483, -28982, -31027, -29626, -27837, -25021, -20965, 
    -18687, -15236, -11398, -6977, -601, 2388, 6584, 10450, 15267, 18942, 
    21692, 25287, 26795, 28497, 31802, 28994, 29334, 30915, 28779, 26369, 
    24462, 20854, 19211, 15108, 11845, 6466, 2907, -3016, -6766, -10279, 
    -15035, -18175, -22863, -25279, -26840, -28878, -28989, -30514, -31042, 
    -29657, -28771, -27973, -24023, -21950, -19587, -14133, -12565, -7120, 
    -1926, 1053, 5195, 11328, 13587, 18329, 22168, 23768, 26503, 28545, 
    29849, 31585, 29524, 30463, 29073, 26586, 25515, 22183, 20164, 15786, 
    12103, 6761, 3308, -1897, -6033, -9467, -14686, -17564, -21718, -23622, 
    -26406, -28210, -28701, -30130, -30388, -31728, -29294, -26394, -26078, 
    -23719, -18483, -14315, -12307, -7530, -4524, 632, 4977, 9807, 13680, 
    18478, 20893, 23806, 26533, 28549, 29895, 30699, 30265, 29694, 29257, 
    26780, 25002, 24175, 19463, 16219, 11549, 8236, 3125, -2024, -5548, 
    -9622, -13563, -17554, -22038, -24610, -26359, -27825, -29134, -30931, 
    -31266, -28758, -30388, -27020, -24858, -22766, -19517, -14615, -12005, 
    -6933, -4402, 648, 6290, 8168, 14016, 16863, 20158, 22691, 26110, 29832, 
    31006, 30612, 30515, 30462, 28294, 29307, 24979, 24429, 19560, 16186, 
    13334, 7709, 4618, -527, -4504, -8804, -12807, -15765, -20551, -22548, 
    -26184, -28907, -28964, -30209, -29851, -30033, -28842, -28579, -26633, 
    -23039, -19080, -17079, -11791, -7514, -4422, 193, 4636, 8743, 12530, 
    16704, 20536, 24672, 25840, 27667, 29316, 31499, 30114, 29886, 30207, 
    26682, 25439, 24420, 19943, 16912, 13202, 8175, 4378, 208, -5635, -8738, 
    -12676, -16411, -19967, -23820, -26199, -27465, -29950, -30655, -31182, 
    -30333, -27941, -27093, -25908, -24569, -20090, -17283, -12921, -8884, 
    -4736, 316, 4349, 8762, 12736, 18172, 19514, 22688, 26565, 26298, 30716, 
    31067, 31072, 31980, 28123, 29001, 26110, 24117, 21088, 15915, 13399, 
    8063, 5577, 1482, -4693, -7600, -13436, -15055, -19917, -23606, -26014, 
    -27759, -31276, -30220, -29647, -30631, -29378, -28543, -26224, -24244, 
    -19512, -16546, -12839, -8383, -5401, 77, 4575, 8327, 11940, 14961, 
    21278, 22367, 25809, 28197, 30056, 29620, 30596, 31561, 30587, 28646, 
    27728, 23880, 20166, 16928, 12806, 9461, 6360, 1209, -3733, -8786, 
    -12857, -16871, -20033, -23913, -25439, -28979, -28252, -29928, -30776, 
    -30122, -29535, -29006, -26492, -24835, -19700, -17090, -14320, -9616, 
    -5560, -2028, 4200, 8177, 12217, 15595, 20754, 22805, 25366, 28684, 
    28704, 28806, 31127, 30731, 31026, 28676, 27021, 23918, 21812, 17947, 
    14051, 8342, 5272, 1864, -3504, -6883, -11970, -16521, -17687, -22928, 
    -25849, -27951, -29008, -30514, -30755, -32348, -29856, -28299, -27221, 
    -25095, -20794, -17735, -13750, -10114, -5072, -1310, 4374, 6976, 11511, 
    15710, 18268, 22085, 24832, 27530, 30252, 31804, 30460, 31539, 31146, 
    29910, 26739, 25235, 21184, 16282, 12652, 9588, 6186, 490, -2163, -7138, 
    -11586, -15455, -19819, -22351, -24290, -26243, -28909, -29569, -31408, 
    -30410, -30199, -28571, -27539, -23928, -21379, -17825, -13182, -10857, 
    -6628, -2006, 2732, 5875, 9791, 16458, 18158, 22355, 24342, 28440, 27948, 
    29435, 30807, 30102, 28864, 29166, 27725, 24217, 23492, 17021, 14827, 
    10418, 5276, 1523, -2247, -6563, -11253, -16368, -18326, -21610, -23603, 
    -28016, -28204, -30810, -30420, -31566, -30480, -27539, -26566, -25041, 
    -21552, -17750, -13465, -10720, -6674, -1759, 2725, 6773, 10807, 15236, 
    17190, 20781, 24901, 26358, 28598, 30486, 29883, 29692, 29069, 30657, 
    28240, 26211, 22193, 19621, 15954, 10561, 6630, 1932, -624, -6608, 
    -10632, -14251, -16462, -22278, -23606, -28658, -28809, -30512, -31441, 
    -31755, -30828, -29716, -27228, -24615, -22619, -18038, -15632, -11152, 
    -8220, -1892, 1047, 6197, 9798, 15356, 17754, 21405, 24316, 25419, 29310, 
    29348, 30942, 31924, 28641, 29636, 28685, 25543, 21420, 19559, 15463, 
    12187, 6293, 3082, -333, -4952, -9430, -15151, -16867, -21325, -24408, 
    -27204, -29601, -29714, -31399, -29501, -30291, -28961, -26948, -26651, 
    -21419, -18892, -16918, -11588, -8860, -2568, -134, 4238, 9831, 13856, 
    17249, 21258, 22385, 25277, 28742, 29542, 29005, 29443, 30127, 28662, 
    28001, 25891, 22951, 19227, 15692, 11621, 6917, 2656, -1513, -5256, 
    -9742, -14589, -17830, -20381, -24403, -25677, -28045, -29401, -29636, 
    -30563, -29925, -28448, -26318, -25762, -22648, -20260, -17022, -11212, 
    -6769, -4311, 1063, 5248, 10466, 14078, 16422, 21254, 23641, 26422, 
    28156, 29820, 31587, 31127, 29673, 28052, 27412, 25168, 22384, 18887, 
    14445, 11921, 8613, 3613, -606, -6044, -9182, -13402, -17853, -19964, 
    -24559, -26920, -28141, -30063, -31742, -29773, -30535, -28074, -28538, 
    -27382, -22499, -18458, -15107, -13116, -7176, -4157, 0, 4418, 9529, 
    14461, 17493, 21014, 24060, 25268, 28092, 31170, 30352, 32415, 31674, 
    29498, 27820, 27143, 24281, 20765, 16469, 11663, 9019, 5140, 254, -5606, 
    -10032, -12681, -16764, -21946, -23486, -25197, -27466, -29790, -30506, 
    -30260, -30890, -29862, -27680, -25715, -23892, -18865, -17001, -11479, 
    -9915, -3962, 167, 4988, 8287, 12369, 15980, 19099, 22573, 26248, 28438, 
    29719, 30578, 29832, 29901, 29451, 28666, 25365, 23782, 20985, 17267, 
    12661, 8726, 4811, -1099, -5436, -7514, -11146, -15420, -18915, -22700, 
    -26370, -28035, -28712, -30152, -30148, -30324, -30212, -28520, -26851, 
    -23042, -19921, -15712, -14211, -9097, -3647, 134, 3875, 8375, 11341, 
    15350, 20468, 22334, 24295, 28027, 28598, 31556, 31146, 28960, 29529, 
    28251, 25453, 22710, 20454, 17498, 11669, 10382, 4115, 2200, -4456, 
    -9623, -12727, -15858, -20941, -22669, -23919, -26264, -29987, -30219, 
    -31095, -29872, -30167, -28019, -27669, -23711, -20958, -17072, -13589, 
    -8822, -4638, -534, 4000, 8217, 12299, 15909, 20174, 21823, 25669, 27628, 
    29879, 29835, 32002, 30265, 30875, 29396, 26125, 23822, 21658, 17476, 
    14914, 9526, 5738, 1588, -3430, -8882, -11299, -16128, -18693, -23218, 
    -23996, -26736, -27724, -31318, -29835, -30015, -28649, -28354, -26349, 
    -24744, -20777, -19282, -13770, -10238, -6032, -1687, 2843, 6750, 12045, 
    14893, 19583, 22934, 23630, 28558, 27962, 29727, 30942, 31165, 29996, 
    29077, 26897, 24566, 23030, 18935, 15202, 8288, 6482, 600, -4040, -8979, 
    -10892, -15316, -18959, -22479, -24346, -27313, -30338, -31659, -29647, 
    -30836, -29795, -29065, -27500, -25578, -22567, -18167, -16001, -8781, 
    -7068, -1546, 3801, 6665, 10990, 15764, 18805, 23031, 24141, 26931, 
    27759, 30035, 32271, 31305, 29635, 28940, 27582, 23957, 22551, 18549, 
    13262, 11069, 5224, 1094, -2618, -7209, -11409, -15165, -18454, -22162, 
    -24785, -26101, -28043, -29884, -30925, -30737, -29397, -29425, -26423, 
    -26416, -21782, -18758, -16004, -9412, -6201, -3916, 1818, 7428, 10670, 
    15660, 18343, 22078, 24444, 26856, 27394, 29706, 30945, 30790, 29739, 
    29802, 27245, 25088, 20867, 18462, 15269, 12009, 8473, 2609, -1841, 
    -6536, -10360, -14414, -18915, -21651, -24588, -26966, -28856, -30344, 
    -30005, -29521, -29039, -27366, -26894, -24985, -21759, -20167, -15441, 
    -11233, -8436, -2559, 1558, 7545, 10802, 13729, 18326, 21485, 24185, 
    25930, 27638, 31081, 30032, 31695, 29613, 27576, 28554, 25483, 21949, 
    18819, 14333, 11071, 6256, 3162, -1562, -4839, -10944, -15281, -17451, 
    -22297, -24225, -26086, -29009, -31346, -30147, -31957, -29338, -28660, 
    -26378, -25454, -22568, -18411, -16359, -12026, -7883, -2987, 2051, 6338, 
    9709, 13147, 19187, 20556, 24406, 27467, 27242, 29016, 32388, 31355, 
    31506, 30132, 28003, 26403, 23609, 19556, 16205, 12196, 7801, 3453, 
    -1753, -4053, -9195, -12942, -16772, -22485, -23707, -26225, -28523, 
    -29473, -29674, -30452, -31446, -29335, -27024, -26452, -23989, -19467, 
    -16149, -13282, -7727, -3912, 2238, 5245, 8171, 14877, 16027, 20202, 
    24092, 26966, 29451, 30655, 29928, 30684, 30116, 30881, 27041, 24184, 
    23008, 17794, 15911, 13156, 8682, 2813, -134, -6220, -8869, -12704, 
    -18442, -20959, -23368, -26195, -27877, -30182, -30039, -30983, -29330, 
    -29701, -27678, -25121, -23117, -19752, -16573, -12108, -7627, -4480, 
    198, 4722, 8888, 14835, 15830, 20344, 24007, 27252, 28599, 29995, 29347, 
    32328, 30778, 30470, 27173, 26340, 23676, 20312, 16656, 12452, 8035, 
    2441, 8, -6116, -7621, -12680, -16611, -20634, -23170, -26380, -27063, 
    -29745, -30758, -30902, -29730, -29410, -28075, -25548, -22185, -20150, 
    -17729, -13045, -9128, -4161, -343, 4569, 9636, 12215, 17232, 18772, 
    22295, 25909, 29262, 28593, 30672, 30518, 30216, 28848, 26518, 26379, 
    24532, 20536, 15197, 13748, 7764, 4260, -985, -5757, -8979, -12211, 
    -15535, -21233, -22512, -26946, -27102, -28800, -30683, -30276, -31797, 
    -28828, -27647, -26292, -23263, -21059, -16415, -13196, -9848, -5145, 
    -1471, 3778, 7591, 13469, 17066, 19244, 23152, 25575, 27974, 28621, 
    30629, 31566, 29864, 28500, 29468, 26708, 23957, 19759, 15896, 12343, 
    9362, 5407, 1775, -4113, -9485, -11067, -16531, -20175, -24415, -24624, 
    -26194, -28853, -31685, -30124, -30548, -28979, -28748, -25897, -23454, 
    -21846, -16601, -13050, -9872, -5423, -1663, 3729, 7059, 12441, 16360, 
    19653, 23689, 26234, 27535, 29293, 31355, 31097, 31200, 29413, 28671, 
    26085, 25350, 20650, 17065, 14208, 10201, 5848, 678, -2865, -7758, 
    -11075, -15081, -19802, -22668, -25491, -28023, -29291, -29225, -29172, 
    -30510, -29999, -28674, -26955, -24156, -20763, -17096, -14255, -10800, 
    -6024, -433, 1268, 7286, 12807, 14232, 19150, 21642, 24806, 27479, 28625, 
    31097, 29678, 30607, 29407, 29289, 25996, 22743, 20289, 18208, 13698, 
    11026, 5763, 825, -2942, -6218, -10445, -15955, -17568, -22548, -23291, 
    -27238, -28775, -30624, -30819, -30702, -30087, -29665, -27033, -25291, 
    -21186, -17179, -13920, -11430, -5107, -1551, 2591, 7269, 11151, 14891, 
    18950, 20682, 25917, 27672, 30572, 30009, 30459, 31219, 29784, 29982, 
    26867, 24805, 20201, 19002, 15502, 11291, 6370, 2016, -3448, -7501, 
    -12203, -15760, -18128, -21174, -24853, -26489, -29039, -29106, -31171, 
    -31488, -30780, -28031, -27580, -25827, -22801, -18826, -15011, -11693, 
    -6132, -1172, 1719, 6193, 12569, 14712, 18762, 21614, 24967, 27546, 
    30281, 31575, 30512, 30988, 28858, 28719, 27629, 23944, 20366, 19748, 
    15276, 11798, 6346, 3554, -1120, -5509, -9784, -15129, -18665, -21400, 
    -25484, -26768, -29471, -30821, -30854, -30247, -31043, -29000, -27797, 
    -24799, -21033, -17780, -13879, -11237, -7108, -3691, 1223, 7277, 10842, 
    14091, 16623, 20883, 23750, 26779, 28012, 29909, 31102, 31607, 30528, 
    28051, 26793, 25172, 22439, 17426, 14787, 10982, 7496, 2753, -1900, 
    -6110, -10033, -13918, -18071, -20934, -23716, -25982, -28017, -29855, 
    -29853, -31135, -29625, -29043, -26722, -24762, -22524, -18394, -15480, 
    -10441, -7798, -3057, 1360, 5581, 8906, 15225, 17956, 20243, 24219, 
    25484, 27033, 29646, 29991, 31438, 29045, 30227, 26868, 25897, 22794, 
    18774, 15185, 12424, 8262, 2659, -1920, -5551, -10045, -12696, -18786, 
    -21371, -22923, -25818, -28383, -30397, -30574, -30067, -29836, -29757, 
    -27791, -25990, -22221, -19858, -16059, -11928, -7702, -3490, 394, 4480, 
    9708, 13548, 18901, 20391, 23702, 27819, 27128, 30341, 30748, 29586, 
    30234, 29851, 28629, 24377, 22553, 19832, 15623, 12394, 8427, 3743, 
    -2003, -4370, -9488, -14747, -17521, -20216, -23720, -25460, -28306, 
    -28551, -29771, -29344, -31217, -28930, -26372, -25078, -21758, -20342, 
    -15463, -10882, -8412, -3727, 267, 4440, 8502, 13975, 16329, 19957, 
    23235, 25658, 27349, 29832, 32134, 29498, 29450, 29382, 28757, 25750, 
    23533, 19994, 17214, 14155, 9421, 4830, 684, -4266, -7848, -12988, 
    -17785, -18955, -22672, -25528, -29674, -29636, -30357, -31382, -29465, 
    -29574, -28859, -25672, -23073, -19740, -16331, -13078, -8673, -5078, 
    105, 4922, 7983, 13599, 15463, 19820, 23758, 24542, 28282, 29040, 30604, 
    32365, 31826, 30837, 28662, 26200, 23713, 21954, 16793, 12600, 8329, 
    5484, -909, -5482, -8001, -12365, -17689, -19934, -23142, -26660, -27769, 
    -29048, -30410, -30976, -30441, -30002, -29539, -26374, -22490, -20922, 
    -16017, -12582, -7709, -4446, -1030, 3849, 9623, 11128, 15622, 19190, 
    23751, 24444, 27992, 30478, 30106, 30020, 29269, 30884, 29211, 25779, 
    23852, 19520, 17689, 13406, 10850, 5964, 1149, -4658, -8599, -11926, 
    -15677, -19854, -21384, -24707, -26246, -28561, -30134, -31388, -29693, 
    -29954, -28730, -26601, -24745, -19812, -16447, -12665, -9040, -5277, 
    -1876, 4351, 8403, 11933, 16840, 20898, 22230, 27244, 27193, 28492, 
    30011, 30413, 29442, 29046, 28859, 27157, 23944, 19915, 16676, 12824, 
    8762, 4744, 1658, -4843, -6680, -12642, -16783, -19281, -22239, -25827, 
    -27345, -29838, -31540, -31755, -29387, -29433, -30033, -27134, -24437, 
    -21231, -18968, -14228, -9228, -5727, -3025, 1624, 6485, 13189, 16324, 
    18714, 21258, 24310, 26180, 30088, 30040, 32047, 31797, 31559, 29075, 
    26091, 23035, 20893, 17652, 15850, 9412, 5271, 2282, -2662, -6568, 
    -12100, -16032, -19057, -22315, -25172, -28410, -28381, -30845, -30535, 
    -32388, -29951, -28349, -27242, -24909, -20241, -19644, -14350, -10424, 
    -6710, -1744, 2296, 6987, 11847, 16034, 19182, 22125, 24376, 27071, 
    30609, 30830, 30981, 30306, 29453, 29557, 26699, 24405, 22367, 17627, 
    15044, 10267, 6690, 1917, -3178, -7893, -9410, -15364, -17184, -22770, 
    -24892, -26674, -29387, -28837, -29448, -31028, -30456, -29481, -28127, 
    -24559, -20882, -18650, -13158, -10106, -6844, -2833, 2532, 7242, 10171, 
    14276, 18228, 21058, 24595, 25887, 27778, 30128, 29295, 31295, 30568, 
    28798, 27062, 24707, 21972, 17489, 15514, 11886, 7685, 4044, -266, -5772, 
    -10600, -13844, -19795, -21227, -25443, -26474, -27127, -30070, -30102, 
    -31313, -31507, -29416, -27143, -25033, -22386, -20452, -15328, -10708, 
    -7607, -2767, 2561, 5190, 9136, 14269, 18147, 19978, 23850, 27438, 29425, 
    28203, 29445, 31879, 28916, 29975, 27701, 24015, 21835, 18676, 14700, 
    10928, 7888, 2243, -2158, -5054, -9226, -13901, -17647, -21661, -25151, 
    -25560, -29542, -30889, -31151, -30978, -30210, -29057, -28035, -24346, 
    -23347, -18903, -14578, -10314, -7293, -3448, 1283, 7244, 11053, 12807, 
    16842, 21241, 23928, 26688, 29624, 30842, 30093, 30983, 29884, 28904, 
    27875, 23703, 23183, 19373, 14717, 12144, 8809, 4059, -1132, -3964, 
    -10213, -14455, -17495, -19501, -24138, -27181, -28882, -29310, -29764, 
    -31082, -31199, -30026, -26426, -26029, -22491, -17819, -15574, -11337, 
    -9093, -3156, 110, 4541, 10055, 11754, 18011, 21879, 24367, 26571, 29076, 
    28527, 29216, 30133, 30278, 28676, 27238, 25795, 22406, 19916, 14786, 
    12667, 6502, 3886, -30, -5460, -9513, -12297, -17610, -20257, -22909, 
    -27360, -29210, -29561, -31424, -30584, -28957, -29001, -28794, -25454, 
    -21882, -20939, -15529, -12170, -8248, -3522, 497, 5093, 9292, 13509, 
    17463, 20959, 22662, 26166, 27752, 29568, 30630, 29904, 30899, 30500, 
    28951, 25998, 22189, 19972, 16768, 13007, 9010, 3919, -401, -3783, -9200, 
    -11723, -16801, -19776, -23374, -26013, -29685, -29619, -30995, -31121, 
    -29468, -30021, -27265, -25795, -22842, -20440, -15401, -12946, -8867, 
    -3352, 979, 5198, 8500, 14015, 16221, 20642, 23683, 25864, 26805, 30513, 
    30571, 29742, 31172, 29898, 26768, 25679, 22723, 21032, 16618, 12036, 
    8621, 5500, 1090, -2605, -9743, -11347, -16172, -19942, -24517, -26851, 
    -27761, -28662, -31250, -30627, -31563, -30083, -29283, -25320, -22345, 
    -18960, -18017, -14017, -10125, -4661, -449, 3117, 8570, 12831, 17547, 
    20903, 23359, 26241, 28033, 30825, 31015, 31204, 29077, 29905, 28548, 
    25869, 24081, 20659, 16734, 13127, 8068, 5785, 249, -4508, -6653, -12766, 
    -15522, -19628, -22450, -24206, -28713, -29178, -28811, -31019, -32074, 
    -30483, -29494, -26532, -23518, -21023, -16922, -12933, -10436, -3580, 
    -550, 2549, 7858, 10986, 15717, 19613, 22970, 26429, 28979, 29548, 29191, 
    30976, 30351, 28492, 26810, 26613, 24238, 21795, 18376, 14283, 11241, 
    3645, 1552, -2891, -8994, -12239, -16056, -19708, -22588, -25285, -26486, 
    -29849, -29758, -30840, -29508, -29217, -28721, -26398, -25232, -21055, 
    -18794, -13631, -10170, -5113, -1080, 3967, 5788, 12292, 15425, 19900, 
    21560, 25886, 27257, 29262, 29918, 30932, 31925, 30815, 29072, 25816, 
    24373, 22152, 17489, 15248, 9550, 7043, 874, -3511, -7838, -10302, 
    -15825, -18854, -23194, -26306, -27793, -28628, -30715, -31981, -30181, 
    -31330, -28196, -26460, -25794, -21051, -17730, -14676, -9025, -5324, 
    -2044, 3233, 5959, 10539, 13747, 17601, 21488, 23753, 28271, 27911, 
    30259, 30174, 32060, 29835, 27416, 27363, 25888, 20600, 17535, 14426, 
    10535, 4918, 744, -3769, -7418, -12200, -15349, -17604, -22703, -24069, 
    -28110, -30202, -29585, -29406, -31495, -30644, -30074, -27908, -25180, 
    -21504, -18606, -15508, -9725, -7050, -1251, 1389, 7108, 11183, 14676, 
    19294, 21817, 23541, 27209, 29560, 28950, 32158, 32276, 29236, 29800, 
    27322, 25048, 21131, 18521, 15029, 11587, 6621, 3729, -3552, -6211, 
    -11284, -14024, -18993, -21705, -24146, -27029, -28654, -29002, -30510, 
    -30965, -30807, -28748, -27124, -25812, -20592, -18193, -15401, -10524, 
    -6947, -4078, 371, 5264, 9818, 14020, 17142, 20944, 23732, 25506, 29416, 
    31450, 29956, 30964, 30881, 28661, 26913, 26505, 20787, 19126, 15207, 
    10105, 7012, 3420, -1033, -5747, -11770, -14781, -18048, -21553, -24286, 
    -26593, -27569, -30543, -30262, -29929, -29907, -29840, -29223, -24097, 
    -21661, -19751, -14830, -11817, -6357, -4562, 2094, 7046, 9001, 12951, 
    17599, 20683, 25390, 25455, 29446, 31199, 31833, 30157, 31462, 29300, 
    27471, 25310, 22372, 18371, 15143, 11229, 7418, 4049, -617, -6264, -9229, 
    -13691, -17003, -21469, -23568, -26257, -29491, -29430, -29590, -29918, 
    -30848, -28859, -27066, -23832, -21697, -19016, -17351, -11572, -7091, 
    -3916, -684, 5585, 9340, 13590, 17218, 20153, 23725, 26276, 28250, 31185, 
    29989, 32078, 30374, 29185, 26878, 25305, 23348, 20666, 15940, 11753, 
    8919, 4653, 15, -4818, -8493, -13364, -17709, -20059, -24268, -26072, 
    -29797, -29150, -28996, -31522, -30831, -29237, -27444, -24836, -23661, 
    -19766, -16407, -12892, -9659, -4262, 966, 4515, 9820, 14113, 16808, 
    18873, 24456, 25529, 27945, 28118, 31002, 31323, 31235, 29809, 27181, 
    25971, 21747, 19005, 16033, 12723, 7071, 4135, -944, -5538, -8990, 
    -13526, -18387, -21202, -22553, -26506, -28497, -29351, -30416, -31736, 
    -28805, -29734, -27175, -25667, -22076, -20764, -17587, -12664, -8085, 
    -4769, 646, 2630, 7629, 13056, 15675, 19411, 22746, 25868, 28885, 29131, 
    31360, 29876, 31272, 28625, 28101, 26268, 21586, 20429, 16866, 12088, 
    9473, 3894, -1350, -5081, -10030, -13729, -16706, -19003, -22983, -24833, 
    -27031, -29789, -31806, -31553, -31460, -29826, -26643, -26827, -22138, 
    -20658, -18655, -13983, -8548, -4151, -949, 3314, 7227, 13185, 15112, 
    19790, 22471, 25767, 27803, 29155, 31398, 30259, 29666, 29939, 27835, 
    26042, 24202, 22413, 18345, 12440, 10100, 4126, 856, -3865, -6826, 
    -12681, -17260, -20219, -22400, -25628, -27440, -28892, -29975, -30410, 
    -30571, -29758, -30201, -26671, -24343, -21426, -17218, -13798, -9619, 
    -5558, -1296, 4037, 7548, 11219, 15545, 20984, 21964, 25302, 29067, 
    28610, 31230, 30146, 29566, 30037, 29208, 26961, 24920, 19868, 17703, 
    12709, 9775, 5489, 1155, -2220, -6466, -11927, -16161, -20472, -21509, 
    -24538, -28170, -28687, -29742, -28916, -31331, -29131, -29584, -27535, 
    -25128, -20651, -18931, -14400, -10204, -6425, 141, 2889, 6195, 10434, 
    15164, 20301, 22588, 23676, 28219, 29214, 30105, 30090, 29903, 30997, 
    27848, 25163, 24801, 21371, 17592, 14915, 8968, 4430, 912, -2868, -7421, 
    -12243, -15315, -17922, -23353, -25576, -26183, -28516, -30264, -30106, 
    -30663, -29853, -28605, -26786, -23854, -21767, -17016, -13970, -10205, 
    -6284, -430, 2643, 7065, 11389, 13873, 19864, 23233, 25980, 28095, 29334, 
    31094, 31048, 30322, 28732, 29022, 26788, 24389, 22157, 18133, 14888, 
    11742, 7484, 1872, -2221, -6757, -10541, -13833, -19610, -22542, -25856, 
    -27323, -28973, -31263, -31472, -30988, -29879, -29481, -27803, -26370, 
    -21468, -18888, -15139, -11646, -7305, -2322, 2707, 6071, 11863, 14834, 
    17058, 22089, 24197, 27243, 28554, 29751, 31420, 29820, 31647, 29009, 
    27978, 24770, 23260, 20174, 13891, 11762, 6201, 2103, -3549, -5897, 
    -10832, -13551, -19165, -20233, -24151, -28028, -28544, -30048, -31084, 
    -31164, -29088, -27401, -28120, -23787, -20939, -18894, -16527, -10585, 
    -7528, -3694, 2234, 5567, 10227, 15797, 17876, 19874, 24358, 25340, 
    29817, 31439, 29431, 30676, 30239, 29010, 27492, 24238, 22967, 18287, 
    16143, 10813, 7953, 3116, -1462, -7138, -10435, -13354, -17735, -22127, 
    -26034, -26659, -28524, -28711, -30300, -29560, -31742, -28933, -27479, 
    -24255, -22009, -20085, -16434, -10894, -6264, -1459, 2747, 6885, 10252, 
    13539, 18633, 20647, 24638, 26183, 29414, 29291, 30865, 32243, 30324, 
    29172, 27127, 26147, 23333, 18612, 16135, 11599, 7949, 4845, -1897, 
    -6772, -9971, -13730, -16261, -21376, -24239, -27570, -28669, -30184, 
    -31149, -31521, -30034, -30059, -28623, -24922, -21851, -19577, -15074, 
    -11293, -8025, -3376, 559, 4344, 9881, 13668, 18323, 20465, 24067, 26584, 
    27872, 30285, 31033, 30028, 31375, 29863, 27799, 26846, 22603, 19227, 
    16572, 11982, 7415, 4013, 193, -4247, -10264, -14015, -16016, -20852, 
    -24234, -26195, -27264, -30862, -30297, -30096, -28896, -29726, -26876, 
    -25233, -23713, -19634, -15347, -12330, -7503, -5610, 95, 4021, 8973, 
    12720, 16865, 20816, 22945, 24233, 28698, 30305, 29313, 29874, 31567, 
    30539, 28999, 24491, 22698, 19232, 16653, 12359, 7960, 3690, -84, -4030, 
    -7755, -12071, -17663, -18998, -23597, -25755, -27466, -29272, -30999, 
    -30008, -30507, -30246, -27446, -27100, -24827, -19835, -16319, -12168, 
    -8074, -3829, -489, 5134, 8757, 12798, 16756, 20194, 22822, 25052, 28859, 
    31446, 29587, 32481, 30426, 30053, 27791, 25449, 24553, 19547, 15442, 
    12804, 9333, 4860, -143, -4359, -9872, -12233, -16940, -21398, -23002, 
    -27205, -26672, -29405, -30270, -31312, -30925, -28471, -28223, -27773, 
    -24219, -19417, -16927, -12596, -7773, -4810, -850, 4243, 8875, 12444, 
    16482, 18793, 22060, 26751, 28201, 29719, 30472, 29107, 30945, 28456, 
    28955, 24923, 22971, 19338, 16667, 13642, 8671, 5293, 1808, -3966, -8087, 
    -12355, -14422, -19816, -24084, -25520, -27738, -28975, -29857, -31009, 
    -30840, -30781, -28323, -26810, -23249, -22060, -16250, -13826, -9036, 
    -3493, -208, 4786, 7827, 10565, 17009, 18823, 22606, 25229, 28690, 29458, 
    30631, 31773, 29596, 30199, 29401, 25995, 24311, 21692, 17509, 13578, 
    8930, 5681, 1837, -3458, -7868, -10780, -16045, -18354, -23888, -25893, 
    -27356, -27605, -30215, -30992, -31233, -29699, -29356, -25763, -22729, 
    -21719, -18186, -13717, -9525, -5288, -1509, 2854, 6813, 11890, 16172, 
    18512, 22639, 24356, 27307, 28079, 29688, 31068, 31096, 29419, 29300, 
    27055, 24820, 21293, 18272, 13181, 9388, 5589, 456, -3308, -6589, -11850, 
    -14701, -17341, -21476, -25451, -26313, -29666, -30800, -30927, -31479, 
    -29543, -29388, -28348, -24446, -20051, -17154, -13267, -10916, -6061, 
    -2493, 1561, 7247, 10500, 16138, 19233, 22384, 25852, 27917, 27579, 
    30620, 31202, 31594, 29671, 29114, 28205, 23464, 22724, 17960, 13971, 
    11169, 6693, 624, -2307, -6964, -10522, -15045, -17150, -23075, -24581, 
    -26616, -30105, -30837, -31329, -29883, -31791, -27119, -25531, -23406, 
    -22917, -19276, -14843, -10688, -7605, -835, 1678, 5866, 9837, 14880, 
    18524, 21605, 24511, 27366, 28060, 29985, 30169, 30547, 30164, 28110, 
    25487, 24560, 23294, 19096, 15112, 10654, 5810, 1403, -2356, -5656, 
    -10522, -14126, -18603, -22445, -25160, -27166, -27985, -28633, -31306, 
    -30529, -30633, -30444, -27789, -25881, -21859, -19349, -15063, -11878, 
    -6401, -3677, 1454, 6822, 11116, 12675, 18196, 22490, 24290, 26381, 
    28529, 29065, 32450, 30409, 30948, 28176, 26044, 24358, 22584, 20382, 
    15422, 11810, 6874, 2753, -2068, -5726, -9930, -15505, -18037, -22550, 
    -25380, -25744, -26883, -31111, -30668, -31171, -30376, -28538, -27840, 
    -25157, -22692, -19103, -15647, -10016, -8105, -4572, 1784, 4151, 10976, 
    14253, 18314, 20380, 24804, 26354, 29156, 30889, 30140, 30041, 29816, 
    29433, 25829, 26306, 21799, 18604, 14908, 12791, 7160, 4036, -587, -6216, 
    -10575, -12794, -18403, -20775, -22830, -27323, -28021, -28819, -30572, 
    -31056, -30308, -28602, -28042, -26340, -24037, -18757, -15324, -11635, 
    -9503, -3715, 1196, 6505, 10288, 12954, 16573, 21207, 22847, 25655, 
    27225, 30968, 32178, 31223, 30411, 29193, 27663, 24736, 22630, 19759, 
    15817, 13425, 6364, 3973, -1877, -5851, -8494, -12529, -17535, -19911, 
    -23888, -27585, -27758, -29753, -28847, -29519, -29492, -28942, -27423, 
    -25050, -21627, -18745, -15836, -12443, -8151, -3368, 59, 5036, 8906, 
    13284, 16844, 21522, 23154, 27123, 28141, 30851, 30897, 31070, 30384, 
    30182, 27705, 26907, 23678, 20544, 17361, 12497, 9340, 3994, -75, -5270, 
    -10115, -12845, -16321, -20179, -22517, -26096, -27225, -29515, -31317, 
    -30878, -30078, -29456, -28663, -25425, -24752, -20023, -16754, -12920, 
    -8612, -5704, -1545, 4936, 9610, 14097, 15917, 19152, 21485, 27568, 
    26803, 29814, 30288, 31470, 30469, 30782, 28652, 26017, 24182, 20458, 
    15797, 14252, 8924, 5279, 1635, -3911, -8158, -13715, -15726, -19527, 
    -22291, -26339, -28857, -30556, -30605, -32336, -31402, -30945, -28046, 
    -25599, -22647, -20949, -16621, -14974, -9752, -5346, -567, 4014, 7998, 
    12691, 14979, 21404, 24119, 26234, 27346, 29679, 30997, 32476, 31400, 
    28381, 29120, 26152, 23367, 19814, 17621, 13055, 9103, 5318, 834, -5156, 
    -8498, -12144, -16221, -20224, -21993, -26541, -27573, -28855, -30097, 
    -31800, -30398, -29097, -27298, -26972, -25242, -20485, -16511, -13217, 
    -8062, -5671, -1860, 3815, 7120, 12280, 15076, 19760, 22193, 24990, 
    27444, 29431, 30413, 31037, 30338, 30011, 30035, 27937, 23180, 21153, 
    19239, 14480, 10736, 5627, 1251, -2530, -7028, -13393, -15766, -20410, 
    -23060, -26506, -27688, -28302, -29541, -30362, -30265, -30322, -28403, 
    -26495, -22757, -21888, -18268, -13989, -9246, -6464, -2308, 2793, 6392, 
    11512, 14035, 18492, 21892, 26102, 27362, 29038, 30036, 30933, 30425, 
    29482, 28891, 25304, 24740, 20444, 19188, 15099, 10446, 5397, 2186, 
    -3319, -5851, -11575, -14110, -19721, -21986, -25247, -27316, -28350, 
    -30552, -31360, -30185, -31131, -28915, -24957, -25458, -21342, -17374, 
    -13999, -11135, -5686, -709, 2558, 5554, 10986, 14553, 18104, 21698, 
    25629, 26871, 28939, 30680, 30804, 32353, 30644, 29036, 27096, 24268, 
    21148, 18208, 14821, 10622, 6298, 995, -2125, -6646, -9637, -13682, 
    -17652, -20689, -24910, -26528, -27708, -30953, -30227, -31087, -29143, 
    -29415, -26077, -24233, -20383, -19634, -14472, -10416, -5566, -2313, 
    2013, 6201, 9544, 14315, 17710, 22173, 23821, 27519, 29021, 31106, 31160, 
    31289, 29369, 29079, 27601, 24109, 20542, 18841, 15154, 11506, 5157, 
    2888, -3510, -6465, -10654, -15149, -20135, -21810, -25471, -26325, 
    -28513, -31257, -32035, -30216, -30634, -29781, -28273, -23554, -23282, 
    -19490, -14402, -11794, -5620, -2481, 717, 5060, 9835, 15057, 18882, 
    21669, 25314, 26637, 29057, 30031, 31186, 30792, 30031, 29270, 27167, 
    25743, 22811, 18693, 15027, 10520, 7507, 3033, -2358, -5673, -11555, 
    -15382, -17503, -20638, -25764, -26115, -29341, -29974, -30642, -29807, 
    -31406, -29856, -28607, -26342, -21299, -17665, -13975, -10408, -5844, 
    -1896, 1733, 6212, 9754, 13657, 17329, 21261, 23302, 26392, 28662, 29607, 
    30860, 30989, 30386, 27695, 27061, 24297, 22481, 18788, 15844, 10859, 
    7622, 3144, -1668, -4713, -10946, -13717, -17315, -20810, -24975, -25598, 
    -28386, -29127, -31076, -30695, -31162, -28626, -29144, -25141, -22117, 
    -19887, -16580, -11697, -8474, -2861, 429, 5623, 8958, 12163, 17452, 
    19484, 24026, 26821, 28706, 30643, 30684, 29859, 31259, 29584, 27713, 
    25855, 22339, 19727, 16336, 12086, 6938, 2333, -1654, -5242, -9642, 
    -12836, -17446, -21365, -22692, -27103, -27185, -30524, -29687, -30294, 
    -30876, -29751, -28245, -24876, -21469, -20521, -15729, -12839, -8535, 
    -4111, -35, 4331, 9066, 13749, 17215, 20168, 22179, 26158, 28349, 29281, 
    30902, 31821, 30163, 28913, 28427, 25424, 23683, 19371, 16654, 13853, 
    8664, 4951, 931, -3991, -7796, -14322, -18511, -19826, -23321, -26781, 
    -26983, -28643, -29711, -30774, -30662, -30053, -27915, -27238, -23835, 
    -19756, -15500, -11926, -8240, -3893, 1053, 3671, 7536, 14279, 15882, 
    20383, 24440, 26479, 27435, 28715, 30245, 30561, 30021, 28418, 28559, 
    25248, 21896, 19694, 16119, 13301, 8009, 4631, 1335, -4582, -8345, 
    -12755, -15420, -19660, -23501, -25692, -27591, -29265, -30161, -30257, 
    -30045, -29895, -27999, -27197, -24746, -21822, -16512, -11767, -8522, 
    -3547, -1002, 3893, 8554, 12839, 15439, 19250, 21977, 25306, 26428, 
    31031, 30001, 32170, 31818, 29939, 28195, 25385, 22924, 19572, 16362, 
    13644, 9159, 4785, 2071, -4578, -7337, -11663, -14668, -20715, -23325, 
    -25850, -26692, -29711, -30722, -31951, -30699, -30434, -28671, -27511, 
    -22743, -20091, -17887, -14459, -8844, -5714, -2275, 2280, 8171, 12043, 
    17605, 18513, 22699, 26093, 27851, 28530, 29864, 29250, 30666, 30131, 
    28344, 27449, 24282, 20705, 16146, 12829, 10638, 5545, 465, -2465, -8075, 
    -10831, -15180, -19885, -22498, -24797, -27413, -28735, -31313, -30486, 
    -31864, -31358, -29509, -26497, -24028, -21545, -17811, -14532, -9423, 
    -5278, 40, 4424, 6158, 12048, 14588, 18711, 20855, 24968, 27466, 29543, 
    31024, 30854, 30838, 29280, 26774, 26166, 24717, 21358, 17419, 13076, 
    9646, 5786, 1019, -3143, -6572, -11540, -14931, -20018, -20865, -26225, 
    -26967, -29116, -30190, -31750, -30151, -31048, -29042, -27674, -24300, 
    -23134, -18417, -15846, -10064, -6063, -2627, 3870, 7662, 11842, 16224, 
    18788, 20550, 24157, 28339, 27424, 29083, 31714, 31120, 29928, 28887, 
    25738, 23693, 21312, 17233, 14404, 9784, 4662, 1991, -624, -6671, -10692, 
    -16081, -17937, -23322, -25796, -27125, -29079, -30306, -30469, -31492, 
    -29179, -28693, -26573, -24094, -21651, -17572, -14053, -9482, -6888, 
    -2097, 2133, 6886, 11981, 14476, 19073, 21852, 25505, 27179, 29290, 
    31754, 31515, 31113, 31113, 28972, 26551, 26188, 20470, 18649, 15432, 
    10805, 6547, 2886, -1986, -6482, -10914, -13121, -18209, -21870, -24683, 
    -25783, -29751, -30613, -31017, -30537, -29805, -29421, -27172, -25194, 
    -22173, -18663, -14485, -10925, -5638, -2148, 990, 7201, 11040, 13510, 
    17957, 21955, 25449, 25478, 27912, 29403, 30346, 31159, 31848, 27896, 
    28905, 25648, 22825, 19739, 15645, 11485, 7974, 1743, -1315, -6689, 
    -9807, -14542, -16309, -20954, -24148, -26455, -27560, -29506, -31799, 
    -29408, -31314, -28852, -27737, -25569, -23644, -19430, -15561, -12752, 
    -7690, -3001, 2065, 5805, 9312, 14582, 17793, 21704, 25053, 26538, 27546, 
    31219, 29508, 31824, 30226, 30869, 28456, 25328, 22446, 19632, 15218, 
    12002, 7448, 3583, -764, -5729, -11040, -12505, -17251, -20471, -24484, 
    -26922, -28479, -28756, -31482, -29716, -30486, -28604, -28518, -26466, 
    -24388, -18845, -15994, -13097, -7607, -3811, 118, 5086, 10121, 14052, 
    18670, 19960, 24017, 26200, 28462, 30894, 29887, 30938, 29810, 29177, 
    26756, 26089, 22018, 20153, 16320, 11956, 6970, 5059, -999, -5190, -8724, 
    -13269, -17776, -20690, -24465, -25827, -27802, -30158, -31850, -30923, 
    -30926, -30465, -26329, -24440, -22273, -20546, -16666, -13063, -8262, 
    -3686, -860, 4081, 8941, 14522, 17507, 21071, 23900, 26407, 28473, 30165, 
    31795, 29863, 29992, 30028, 27674, 25383, 23681, 19236, 18075, 11777, 
    7257, 3895, 89, -4032, -7258, -13660, -16237, -19874, -23209, -25883, 
    -27302, -30711, -29452, -31104, -28648, -29130, -27106, -27190, -23145, 
    -19281, -17148, -12645, -7396, -3169, -1168, 3040, 9286, 12138, 16382, 
    20514, 23105, 26888, 27871, 28786, 30424, 31496, 29473, 29517, 27520, 
    25474, 23280, 19365, 16889, 13642, 10238, 3929, 415, -4931, -8631, 
    -11071, -17136, -20144, -22527, -23950, -27632, -28019, -31081, -32099, 
    -29246, -28777, -27843, -25178, -24467, -18925, -16601, -12964, -9938, 
    -4306, -1919, 3632, 8923, 12602, 16804, 19169, 23020, 24153, 28050, 
    29604, 30250, 31984, 29252, 29862, 27986, 25610, 23563, 21947, 15998, 
    12213, 9433, 4148, -136, -3649, -7947, -12029, -16720, -20240, -23945, 
    -24944, -27039, -30042, -30863, -31542, -30576, -29016, -28197, -25930, 
    -24726, -21843, -17084, -15086, -9704, -5335, -111, 4755, 7002, 11670, 
    15376, 19632, 22030, 25529, 27689, 27566, 29818, 29397, 29296, 28881, 
    29185, 27329, 23554, 21197, 17043, 14017, 8954, 4704, 86, -4140, -8932, 
    -12065, -16263, -20431, -22292, -25097, -28319, -28426, -30586, -30920, 
    -31179, -30779, -28937, -26636, -23590, -20675, -17667, -15468, -10454, 
    -7538, 283, 3726, 6795, 10184, 16544, 18154, 22626, 23850, 26232, 29361, 
    29338, 31968, 30573, 30413, 28027, 27599, 23024, 20850, 16985, 15542, 
    10966, 6634, 1945, -3044, -6822, -11061, -14464, -20120, -21193, -24901, 
    -26852, -28667, -29423, -32462, -31419, -29059, -28959, -26088, -24517, 
    -21702, -18725, -13523, -10521, -5082, -1892, 2771, 6308, 11109, 13697, 
    17474, 22503, 24137, 26879, 27859, 31972, 30817, 30736, 30900, 29703, 
    27054, 24485, 23183, 18139, 15813, 10411, 7196, 458, -1882, -6765, -9664, 
    -13921, -17904, -21803, -25010, -26308, -28301, -29682, -30685, -31224, 
    -29483, -28616, -27409, -26163, -22052, -18931, -13850, -11225, -6442, 
    -3448, 1465, 7825, 12185, 14518, 19720, 22645, 25094, 27428, 28548, 
    29108, 30539, 31020, 30765, 29556, 26035, 25027, 23388, 18300, 14902, 
    10632, 6380, 2630, -2241, -5772, -10046, -14505, -17921, -21763, -24586, 
    -27642, -28603, -29448, -31627, -32194, -30388, -29634, -27644, -24017, 
    -20440, -18605, -15365, -10248, -5781, -3578, 2275, 5593, 9787, 15308, 
    16899, 21335, 23423, 26188, 28847, 29814, 30669, 30958, 29753, 29416, 
    27972, 25123, 22879, 19793, 15824, 11299, 7111, 2002, -1447, -6230, 
    -11347, -14977, -19222, -20476, -24029, -26343, -29291, -29301, -31760, 
    -30479, -28682, -27750, -27281, -24168, -22560, -19613, -14479, -11028, 
    -7291, -1341, 1997, 6070, 10049, 13693, 17806, 21265, 23502, 25446, 
    29951, 29582, 30030, 30414, 31491, 30162, 28625, 25320, 22694, 18632, 
    16216, 11410, 7180, 3282, -2330, -6608, -9468, -13166, -17256, -20962, 
    -24269, -25730, -29540, -29821, -30423, -29582, -32049, -29160, -26659, 
    -24521, -21688, -19975, -16586, -11268, -7259, -3374, 228, 4908, 8404, 
    13078, 18115, 20642, 23257, 26690, 28774, 29110, 30560, 31101, 32036, 
    29600, 26262, 26305, 22233, 20370, 17064, 13730, 8194, 3697, -150, -6235, 
    -9026, -14381, -17537, -20560, -22714, -25435, -29491, -29560, -29142, 
    -30320, -30809, -30519, -28682, -25656, -22536, -20556, -16898, -13299, 
    -7718, -4859, -444, 4295, 9465, 12999, 18529, 19316, 24792, 27288, 28840, 
    29278, 30964, 29871, 31237, 29586, 27426, 26548, 23340, 18570, 17288, 
    13214, 8480, 3040, -1102, -4740, -8572, -13128, -16728, -19597, -23221, 
    -25976, -26403, -29343, -31428, -30992, -30515, -30528, -28416, -26627, 
    -22849, -20653, -16778, -11626, -9202, -5962, -561, 4508, 9491, 12598, 
    17224, 20567, 23178, 26385, 27356, 29518, 29575, 30929, 30028, 29060, 
    26991, 27252, 24190, 19408, 17593, 12136, 7168, 5444, 1432, -3915, -7701, 
    -12218, -15328, -18877, -23297, -24031, -28796, -29280, -31411, -31918, 
    -30625, -28396, -28439, -25119, -22660, -19841, -17228, -12036, -7879, 
    -3517, -671, 4739, 9456, 11682, 15386, 18796, 21950, 24497, 27073, 29592, 
    30621, 30356, 31103, 30198, 26553, 25119, 24336, 21101, 18001, 13365, 
    9744, 5130, -336, -4238, -8768, -13221, -15283, -19611, -23117, -25753, 
    -28311, -30138, -30154, -30753, -30859, -30569, -27474, -25878, -24352, 
    -20326, -16732, -12326, -8715, -6468, -660, 3397, 8202, 13220, 14482, 
    19752, 22865, 26510, 28223, 28950, 30584, 31259, 29398, 30459, 29059, 
    27997, 23457, 22000, 18768, 13164, 9770, 6636, 1910, -3838, -7492, 
    -11288, -14203, -19937, -21438, -25533, -26476, -29386, -29146, -29928, 
    -30277, -30738, -28936, -26308, -25406, -20082, -17396, -14633, -9972, 
    -5212, -1489, 3778, 8709, 11753, 15020, 19483, 22929, 24734, 27744, 
    29459, 31269, 31205, 31241, 29719, 29037, 27240, 23497, 20423, 16941, 
    12914, 9011, 5705, 2471, -1802, -7312, -11832, -15614, -17761, -21728, 
    -24166, -26983, -27434, -30101, -31004, -30722, -29189, -28580, -25865, 
    -25258, -21993, -17935, -14893, -9567, -7460, -1596, 1754, 6392, 10491, 
    14783, 17770, 20683, 26203, 27739, 29904, 29071, 30562, 30249, 31069, 
    27617, 25983, 24482, 21779, 17966, 14818, 9851, 6614, 1479, -3943, -7047, 
    -10780, -14416, -19911, -23213, -24144, -26505, -28531, -29423, -31426, 
    -31037, -29334, -29866, -26222, -24848, -20174, -18823, -14195, -11922, 
    -6583, -3495, 2117, 6052, 10687, 14383, 19416, 21976, 25050, 25950, 
    27765, 29016, 30629, 31341, 29472, 29564, 26082, 23763, 21874, 19626, 
    15178, 11133, 7915, 2918, -1823, -6538, -10290, -13950, -16792, -22145, 
    -25461, -27367, -28533, -30626, -31495, -29545, -28884, -28685, -26095, 
    -24730, -21763, -20157, -15058, -11978, -6806, -1453, 3364, 5329, 10254, 
    14538, 17561, 21944, 24929, 27146, 30221, 31113, 31285, 31489, 31040, 
    28171, 28210, 26395, 22787, 18777, 14682, 11250, 7121, 4372, -862, -6927, 
    -9682, -12426, -17795, -21317, -23831, -27383, -28444, -30061, -30166, 
    -30883, -29008, -29687, -28204, -25603, -22559, -19991, -14306, -12726, 
    -6124, -2645, 1398, 4834, 9684, 12872, 17323, 21493, 24039, 26778, 27744, 
    31770, 30086, 31110, 30989, 30483, 27538, 25914, 22979, 19582, 16517, 
    10789, 8805, 1844, -346, -3659, -10460, -15122, -17184, -20635, -24940, 
    -25750, -28986, -28378, -29096, -31969, -30364, -30053, -27314, -25434, 
    -21989, -19011, -15877, -12141, -6915, -4135, 2501, 4242, 9684, 13826, 
    18141, 19959, 22966, 27228, 29403, 30539, 30609, 31324, 30003, 29559, 
    28406, 25426, 24417, 17893, 16265, 10777, 8882, 3794, -1110, -5239, 
    -10177, -12079, -16879, -19837, -22278, -25508, -29558, -28863, -31361, 
    -31764, -31578, -29014, -27868, -24856, -23047, -19843, -16889, -13910, 
    -7598, -5318, 795, 3685, 10278, 12827, 17001, 18941, 22325, 26342, 27720, 
    28632, 30863, 30769, 30659, 28708, 27375, 27105, 23655, 18242, 16531, 
    12397, 7565, 3884, -136, -5824, -8412, -12644, -18597, -19752, -24009, 
    -26788, -27666, -30442, -28979, -29856, -30127, -30080, -29107, -25268, 
    -22984, -21025, -15590, -13390, -8401, -5264, -39, 4687, 7492, 12996, 
    15081, 19841, 23828, 24905, 27161, 28856, 28714, 31623, 29491, 30286, 
    26933, 27061, 21885, 21138, 17810, 14262, 8218, 5720, 787, -2994, -9384, 
    -12467, -16484, -20167, -22063, -26374, -28569, -28948, -29813, -31366, 
    -29557, -30149, -28148, -25479, -21977, -21188, -17835, -13205, -9819, 
    -4509, -551, 2838, 7030, 12238, 16127, 20898, 23044, 25884, 27447, 29258, 
    30697, 29594, 29938, 29800, 27281, 25244, 24753, 21571, 16602, 15051, 
    9908, 6281, 1463, -2424, -9477, -11540, -15509, -20096, -23870, -25516, 
    -26269, -28571, -30520, -30962, -31631, -28553, -27442, -24665, -22561, 
    -21767, -16847, -14054, -9619, -5297, -2285, 3272, 8313, 11202, 16556, 
    19566, 21158, 25376, 27777, 27949, 31209, 30639, 31488, 28998, 27401, 
    27100, 24222, 20633, 16673, 13702, 9178, 6077, 1406, -1650, -8588, 
    -11316, -17299, -20522, -22405, -26582, -27695, -28554, -30811, -32333, 
    -30915, -28801, -27162, -27768, -23734, -22439, -18166, -13792, -10060, 
    -4612, -1127, 4617, 7471, 12999, 16479, 18304, 22607, 24480, 28583, 
    29361, 30075, 32217, 31943, 30954, 29503, 25306, 24652, 21090, 18440, 
    14956, 9119, 5211, 1378, -3475, -6402, -12326, -14224, -17861, -21146, 
    -24353, -28847, -27852, -30705, -31234, -31208, -31081, -27804, -26098, 
    -23300, -20917, -18444, -14754, -10045, -7089, -607, 1839, 7629, 10774, 
    14662, 18217, 22528, 25115, 27003, 28648, 30184, 31256, 31134, 30800, 
    29374, 27670, 25606, 20545, 19526, 14973, 10440, 6752, 2498, -711, -6930, 
    -10341, -15078, -17390, -22563, -23075, -26376, -28330, -30204, -30111, 
    -31393, -31110, -27437, -27022, -24601, -21017, -17738, -14090, -9404, 
    -5380, -2346, 2251, 5365, 9748, 14687, 18030, 20920, 25362, 27397, 30616, 
    28836, 29697, 30277, 29274, 27637, 28161, 25588, 21586, 18737, 15624, 
    11808, 7926, 973, -2215, -6053, -10508, -14882, -19911, -21008, -24847, 
    -27704, -28738, -29471, -31819, -31178, -29153, -29157, -27769, -24297, 
    -21770, -18733, -15957, -11750, -7652, -880, 2135, 5863, 11886, 13121, 
    18427, 22720, 24028, 26127, 29243, 29956, 31771, 30822, 30256, 30796, 
    26070, 25270, 23974, 17576, 16919, 9663, 6390, 3717, -3055, -6742, 
    -10871, -13747, -18656, -21341, -24313, -26659, -28896, -29469, -29967, 
    -29570, -29831, -29594, -28593, -25884, -22574, -18624, -15043, -12244, 
    -7269, -2278, 1758, 6457, 9771, 12455, 18106, 21849, 22793, 26928, 27568, 
    30559, 31091, 30898, 30023, 30417, 27169, 24409, 22160, 19370, 16707, 
    13126, 7970, 2681, -1808, -3681, -9711, -12924, -18026, -19183, -25242, 
    -26235, -28504, -31169, -30808, -31594, -28809, -29286, -28940, -26509, 
    -22987, -19020, -15563, -11134, -7372, -2461, 468, 4981, 9145, 12211, 
    17145, 21694, 23979, 26656, 27928, 30068, 30261, 30962, 29360, 30421, 
    28851, 26059, 21773, 18148, 17687, 13698, 6684, 3101, -846, -5297, -9475, 
    -13261, -17849, -20504, -24524, -26853, -28424, -29390, -30954, -30247, 
    -31057, -29921, -27970, -25640, -23027, -18809, -15757, -12206, -9019, 
    -4851, 1028, 5653, 8232, 13138, 15976, 20119, 21995, 25806, 27534, 29419, 
    30901, 31218, 29619, 29173, 28099, 26675, 22547, 20112, 16422, 12803, 
    8998, 4635, -1278, -3804, -9530, -12215, -15621, -18969, -23884, -26778, 
    -26581, -28524, -30520, -31690, -30729, -30146, -27527, -26439, -21992, 
    -21132, -18131, -13982, -9531, -5474, -151, 3142, 7628, 13153, 17774, 
    19259, 23460, 24948, 29118, 29665, 30898, 32411, 32193, 30250, 28979, 
    27133, 24130, 21844, 17142, 11880, 8992, 5321, -327, -4034, -9134, 
    -11065, -16980, -20390, -24586, -24947, -27976, -29577, -31246, -30377, 
    -30409, -29603, -27796, -25981, -23613, -19467, -16889, -13033, -9097, 
    -5774, 53, 4982, 8091, 12531, 16757, 19282, 22135, 24559, 27768, 30122, 
    30940, 32263, 31668, 29407, 28250, 25756, 23592, 19124, 17857, 13690, 
    7761, 5057, 1106, -2230, -8924, -12888, -15606, -19090, -22614, -24305, 
    -27972, -29366, -31183, -31350, -29731, -29594, -29311, -27306, -24200, 
    -19164, -16900, -13614, -8150, -4496, -1188, 4915, 7813, 12752, 15124, 
    19435, 23899, 26313, 28379, 27964, 30826, 31133, 29863, 30182, 29654, 
    26402, 24131, 21098, 17355, 15351, 8983, 6644, 2019, -4184, -7096, 
    -11321, -14388, -19439, -21839, -25886, -27140, -27975, -29606, -30228, 
    -30049, -30341, -29587, -24795, -24577, -20607, -18221, -14494, -11053, 
    -5653, -564, 4369, 8934, 12943, 14295, 18602, 22649, 26112, 25674, 28967, 
    31106, 31371, 29963, 29902, 28578, 26647, 23856, 21202, 17823, 14473, 
    10145, 6629, 551, -3064, -5744, -10870, -14064, -19028, -22404, -25357, 
    -27204, -28924, -30453, -30621, -29851, -28697, -28029, -26903, -25045, 
    -22305, -18562, -15653, -10839, -7499, -322, 2309, 8022, 11657, 15320, 
    19277, 22370, 24122, 26525, 28652, 30379, 30338, 32085, 30436, 29235, 
    26839, 23507, 22023, 19216, 14825, 10734, 5105, 2431, -2406, -8004, 
    -10819, -15925, -19521, -21254, -23605, -27415, -28158, -30723, -30951, 
    -30412, -29999, -29375, -26944, -24680, -22511, -18184, -13854, -11367, 
    -5620, -1033, 2125, 7449, 10094, 14967, 19368, 21778, 24606, 27058, 
    27909, 31797, 30458, 32285, 29041, 28364, 27018, 23992, 20788, 18974, 
    15976, 10273, 5305, 3690, -2683, -5948, -10977, -15316, -18555, -20925, 
    -24251, -27289, -28786, -30705, -31160, -30237, -29275, -28202, -26825, 
    -25038, -23268, -19471, -14217, -13034, -6216, -2610, 2480, 6840, 10974, 
    14909, 19085, 21807, 23612, 26218, 28690, 29665, 31258, 30743, 30102, 
    27561, 27246, 25352, 21589, 19012, 14088, 11657, 6857, 3973, -9, -5902, 
    -10152, -13087, -17694, -21334, -23852, -27854, -27172, -29182, -30221, 
    -29730, -29875, -28879, -26268, -26548, -23308, -19189, -15088, -10627, 
    -6838, -1912, 1263, 5694, 11079, 14855, 17608, 20944, 23376, 27179, 
    29236, 30526, 30677, 29801, 29174, 29588, 29364, 25276, 21869, 18643, 
    15841, 10431, 6362, 3822, -891, -5641, -10916, -13943, -17234, -21769, 
    -23969, -27574, -28632, -30760, -31873, -30504, -31491, -29106, -28095, 
    -25400, -23062, -18747, -14762, -13063, -6756, -4464, 1014, 5542, 8854, 
    13017, 17055, 19814, 24875, 26612, 28524, 29061, 29742, 29521, 29573, 
    28380, 28580, 26825, 23654, 20588, 14949, 12713, 9130, 3418, -525, -5140, 
    -9347, -13620, -17365, -21416, -22342, -26516, -28668, -30359, -31451, 
    -31306, -30329, -29184, -26480, -24526, -24339, -19372, -16750, -11102, 
    -8091, -3608, 258, 3808, 7649, 13821, 18182, 19412, 23771, 24846, 28280, 
    30166, 30954, 30578, 31281, 29632, 27869, 26224, 22945, 20989, 16766, 
    11836, 7385, 2773, 1487, -4177, -8542, -11793, -15883, -20377, -24000, 
    -25191, -27697, -31243, -30366, -30238, -31417, -30120, -28743, -25624, 
    -22731, -19738, -16099, -13606, -7731, -4831, -108, 4705, 8748, 13776, 
    17541, 20830, 23357, 25804, 28686, 27751, 30345, 30796, 29077, 30120, 
    26647, 25473, 23893, 20281, 17719, 13069, 8522, 5334, 484, -4337, -7374, 
    -11889, -16151, -19232, -23684, -25806, -28798, -28549, -31663, -31376, 
    -30306, -28322, -29031, -25566, -23808, -19887, -17305, -12359, -9160, 
    -5905, -626, 4377, 9740, 12120, 17770, 18647, 23705, 24836, 27487, 27788, 
    30420, 30936, 31564, 29549, 28356, 26940, 23316, 19992, 17278, 13174, 
    8467, 5545, 1163, -3690, -9157, -13599, -16081, -21028, -21809, -26242, 
    -26220, -28267, -32177, -32412, -30258, -30229, -29139, -26882, -22878, 
    -19823, -17692, -13434, -9495, -4695, 203, 4682, 6301, 13198, 15991, 
    21049, 23935, 25178, 28327, 30042, 29320, 30281, 31115, 30266, 28161, 
    27497, 23899, 21007, 17807, 12509, 11180, 7027, 389, -3662, -7488, 
    -11709, -17050, -18203, -21474, -24222, -27402, -29809, -30706, -30291, 
    -30733, -28547, -28721, -25427, -24098, -20525, -18536, -14674, -10355, 
    -5525, -807, 3212, 7085, 12818, 17023, 20871, 23974, 26733, 27216, 28748, 
    30840, 29511, 31653, 30654, 29310, 27687, 23581, 21318, 18061, 13035, 
    10763, 5269, 649, -2756, -7539, -10963, -15808, -18870, -22069, -25872, 
    -28857, -30424, -30857, -31225, -29997, -29495, -29576, -27656, -23164, 
    -21574, -17209, -14698, -9763, -6594, -1251, 4151, 7323, 11326, 14981, 
    18635, 21976, 24085, 25723, 28361, 28723, 31127, 31225, 29713, 29832, 
    26845, 23891, 21092, 17885, 15836, 9983, 6791, 3557, -2421, -7038, 
    -10315, -14354, -17229, -23080, -25586, -25565, -28150, -30772, -32017, 
    -30144, -30028, -28779, -25671, -23495, -21181, -19234, -14660, -10082, 
    -7305, -2770, 1488, 6630, 10630, 15222, 17880, 22895, 25401, 26199, 
    29669, 31270, 29706, 29377, 31128, 28214, 27402, 24187, 21415, 18538, 
    14280, 11135, 6990, 2892, -1763, -6881, -11002, -14778, -18866, -22564, 
    -25275, -26694, -29160, -28870, -31055, -30947, -30504, -29774, -27128, 
    -25722, -22564, -17828, -14658, -10906, -6369, -1750, 2534, 4952, 10776, 
    14985, 18088, 23255, 24204, 26507, 29006, 29108, 30795, 30132, 29389, 
    28571, 27084, 25143, 22529, 18632, 15837, 12216, 6356, 2411, -498, -4741, 
    -11477, -14541, -17982, -19986, -23001, -27090, -28368, -30091, -30051, 
    -30026, -30362, -28699, -27354, -25425, -21353, -20527, -14492, -12128, 
    -6220, -1870, 2354, 5804, 9882, 14641, 18746, 20698, 25081, 27871, 28663, 
    30488, 30457, 30904, 30389, 29796, 28088, 25901, 23564, 19316, 16760, 
    12360, 8739, 4010, -461, -4707, -8672, -13957, -17821, -21484, -23445, 
    -25917, -29385, -31254, -30433, -29329, -30110, -28396, -28586, -24951, 
    -22650, -19975, -16877, -11690, -8213, -3835, 499, 5408, 9451, 12913, 
    17133, 21117, 22259, 26689, 27365, 30019, 31265, 30340, 30731, 29758, 
    26346, 24639, 23689, 19238, 15170, 12864, 7459, 5135, -1761, -6034, 
    -9468, -14402, -16647, -20361, -23644, -26336, -28067, -28259, -30256, 
    -30445, -29914, -29591, -28592, -26306, -21623, -19580, -15589, -11573, 
    -8280, -3348, -260, 4674, 9462, 13270, 17253, 20007, 24334, 27248, 29695, 
    31355, 30592, 29858, 29582, 29031, 27516, 26415, 24752, 20713, 15855, 
    13894, 7842, 3474, 569, -4042, -9592, -13141, -15551, -20817, -24443, 
    -25950, -27600, -29614, -31265, -30392, -30614, -30339, -27285, -26455, 
    -23490, -18882, -17121, -12618, -8648, -5113, 436, 5150, 8804, 12327, 
    16915, 20289, 24106, 26730, 27837, 30480, 31743, 30801, 30335, 30232, 
    27510, 25277, 23694, 19823, 17118, 14529, 8471, 5048, 15, -5101, -9957, 
    -12234, -17039, -19409, -23008, -25238, -28843, -27706, -30946, -31507, 
    -31338, -29820, -27969, -26727, -23146, -20755, -16199, -13734, -8653, 
    -4331, -1702, 2538, 9129, 13066, 17657, 20483, 22342, 26958, 27516, 
    29656, 31275, 31120, 30113, 31060, 27495, 26667, 23928, 19375, 16557, 
    14311, 11114, 6554, 402, -5164, -8183, -12396, -16342, -20041, -21381, 
    -24798, -26966, -30775, -28631, -30437, -31496, -30701, -29383, -27140, 
    -24167, -19667, -16473, -13503, -9638, -3589, -835, 3038, 8480, 10307, 
    16662, 19875, 23839, 24261, 26826, 29472, 29155, 31272, 30167, 30438, 
    28995, 26637, 22900, 19987, 16362, 14298, 10696, 6370, 288, -1860, -6196, 
    -13165, -16510, -20276, -23847, -25036, -26072, -27381, -30166, -30931, 
    -29365, -30325, -27926, -27069, -23297, -21534, -18666, -14255, -10632, 
    -5033, -1685, 2301, 8057, 10724, 15731, 19330, 21350, 26071, 27593, 
    28185, 28713, 31878, 30254, 30293, 28511, 25493, 24438, 22348, 18420, 
    13723, 10095, 5364, 2157, -3151, -6616, -11597, -14866, -17580, -21195, 
    -24388, -27098, -29083, -29736, -29928, -30879, -29843, -28144, -26375, 
    -24591, -21286, -16969, -12984, -10332, -6895, 89, 2746, 6817, 11544, 
    16108, 19667, 21771, 24280, 26836, 30313, 30284, 30867, 30274, 31024, 
    29118, 27414, 25337, 23172, 18908, 13970, 11089, 7205, 3630, -1504, 
    -5758, -11193, -15188, -19942, -22095, -23852, -25915, -28088, -29098, 
    -31322, -29760, -30272, -28456, -27028, -24887, -21744, -17303, -14160, 
    -11529, -6311, -1826, 3188, 5324, 9832, 14807, 19540, 21320, 24468, 
    27155, 29451, 30187, 29888, 31458, 30340, 28288, 27879, 24798, 22312, 
    19926, 16210, 10681, 6550, 3734, -2972, -6555, -9912, -15126, -18089, 
    -22781, -24253, -27467, -29251, -30101, -31069, -30873, -30950, -28713, 
    -27453, -25017, -21882, -19160, -15803, -12404, -6553, -3807, 1596, 7153, 
    9397, 14038, 18689, 21034, 24106, 25286, 29484, 28941, 30485, 31208, 
    29442, 28521, 27839, 25582, 23561, 19237, 14689, 12459, 7809, 2861, 
    -2333, -4761, -10065, -13534, -18468, -21919, -23973, -27347, -28123, 
    -31571, -29988, -29398, -30439, -28558, -29002, -24029, -21125, -19272, 
    -15482, -11916, -7227, -3247, 1226, 6219, 9677, 14594, 16778, 20410, 
    23328, 25398, 28391, 29276, 29802, 29130, 30881, 28087, 26022, 24996, 
    23321, 20919, 14765, 12228, 6526, 4165, 456, -6725, -9233, -14410, 
    -18368, -20401, -23001, -26915, -28376, -28626, -31488, -31258, -29843, 
    -30135, -27386, -25548, -24132, -19693, -16789, -11799, -6634, -4212, 
    756, 4709, 9704, 14602, 17627, 20282, 23555, 26670, 28766, 29770, 29408, 
    30630, 30155, 28730, 28232, 24788, 24035, 20244, 15505, 12288, 7183, 
    2848, -1106, -4900, -9200, -11872, -16555, -19691, -23597, -25554, 
    -28610, -29975, -30097, -29381, -30794, -29635, -25955, -25191, -22741, 
    -18839, -16889, -11249, -8479, -4119, 1391, 5254, 9641, 13605, 17365, 
    21302, 23672, 25913, 28416, 29666, 30027, 30596, 32048, 29321, 28967, 
    25046, 23811, 19195, 15096, 13871, 9435, 4074, -578, -4372, -9784, 
    -12552, -16586, -20671, -23644, -25108, -27120, -29045, -29582, -30936, 
    -30028, -30707, -28090, -25666, -23101, -20533, -17846, -13785, -9668, 
    -4215, -95, 4573, 9880, 12263, 15436, 20021, 23514, 25540, 27967, 29302, 
    31615, 31569, 31512, 28729, 27533, 25352, 23069, 20098, 17730, 12948, 
    9393, 3500, -337, -5171, -7078, -13782, -15071, -19050, -22171, -25051, 
    -27185, -30038, -30493, -30669, -31947, -29186, -28142, -27111, -22763, 
    -20201, -17091, -13208, -7994, -5029, -1333, 4121, 9667, 11595, 17371, 
    20015, 24906, 25510, 28273, 30078, 29061, 30338, 31010, 30142, 28110, 
    25473, 24849, 20718, 16675, 13071, 10152, 6175, 1111, -4496, -9638, 
    -13355, -15692, -20726, -21458, -25948, -29211, -29731, -29851, -29399, 
    -30559, -29428, -28114, -27618, -23240, -20708, -17768, -13056, -10324, 
    -4207, -350, 2741, 7176, 13648, 15641, 21143, 22513, 26432, 27334, 30036, 
    30724, 29304, 30125, 29360, 29629, 25562, 24930, 20527, 17663, 14396, 
    8502, 6086, -12, -3328, -6593, -12005, -16493, -18752, -21857, -25595, 
    -27244, -28965, -31021, -31647, -28841, -30022, -27631, -26199, -23602, 
    -21469, -18235, -13561, -8235, -6537, -2051, 2472, 6869, 11983, 14782, 
    19998, 23353, 26369, 26439, 28660, 29854, 29895, 30260, 29818, 28770, 
    25853, 24786, 22602, 17116, 13874, 10316, 6039, 2849, -3803, -6183, 
    -10527, -15149, -19367, -22936, -25409, -27369, -29026, -30768, -30121, 
    -31375, -29411, -29932, -26223, -24302, -21655, -19506, -14592, -10479, 
    -5282, -1872, 2160, 6950, 10828, 15175, 17635, 21114, 24915, 26112, 
    27334, 29914, 31281, 31067, 29902, 30230, 27853, 24615, 21444, 16784, 
    14677, 10448, 5947, 929, -1238, -6786, -11293, -14717, -18012, -21210, 
    -25584, -27711, -28549, -30110, -31527, -29696, -30082, -28920, -27701, 
    -25636, -21936, -17648, -15217, -9882, -6756, -1000, 347, 5738, 10684, 
    15800, 19022, 22475, 24859, 27414, 29283, 30584, 30593, 30291, 29221, 
    27370, 25290, 23649, 21380, 18491, 13778, 11044, 6187, 2268, -1907, 
    -7283, -10507, -14337, -18538, -20029, -24672, -26132, -28654, -30112, 
    -30361, -30879, -31555, -29739, -25870, -24746, -22837, -18039, -15702, 
    -10955, -6812, -2667, 1541, 5651, 10964, 14567, 18450, 20450, 23629, 
    26903, 27388, 28796, 30394, 30874, 30506, 29015, 27647, 23886, 23406, 
    18361, 16224, 12135, 6583, 3140, -2444, -6255, -10415, -14002, -17974, 
    -20519, -25454, -26464, -28866, -30110, -29865, -30259, -29709, -29013, 
    -27743, -24789, -21610, -19011, -16083, -11349, -6682, -3069, 2551, 5008, 
    10190, 13960, 19370, 19735, 23692, 26683, 28431, 29024, 32082, 30113, 
    31306, 29399, 26813, 25544, 23199, 20039, 15904, 11471, 6847, 3656, -815, 
    -3601, -10596, -14008, -16996, -20764, -23803, -25821, -27401, -28369, 
    -30390, -31270, -30176, -28625, -26430, -25131, -23218, -19314, -15252, 
    -11029, -7909, -2237, 1689, 4915, 9581, 14564, 16893, 20757, 23047, 
    26447, 28275, 29745, 30734, 31632, 30742, 30118, 27429, 25924, 24194, 
    18215, 16639, 13587, 8479, 3480, -16, -4603, -9463, -12932, -17324, 
    -21330, -23315, -27615, -29722, -30986, -31898, -32748, -31159, -28594, 
    -28369, -25649, -22654, -20213, -16349, -12175, -7785, -3712, -308, 3990, 
    8403, 11988, 16667, 20705, 22688, 24789, 29300, 28867, 28925, 29667, 
    29948, 30473, 28116, 25556, 22942, 18650, 15857, 13124, 8399, 4817, -576, 
    -5024, -10141, -13864, -17611, -21540, -23204, -27896, -28404, -30199, 
    -31066, -30295, -30018, -30154, -28606, -25686, -22708, -20323, -15127, 
    -13781, -8868, -3046, 153, 4273, 8536, 12713, 16377, 19936, 21966, 25814, 
    26275, 30598, 30588, 29797, 30081, 29013, 27518, 26095, 23186, 20746, 
    16943, 12613, 9596, 5200, 597, -3906, -9346, -11708, -15698, -20126, 
    -22233, -25468, -28225, -29821, -30579, -31771, -30362, -29606, -29296, 
    -25429, -25030, -20634, -16061, -12547, -9560, -5957, -224, 4989, 6892, 
    12571, 15911, 20102, 23142, 25880, 28659, 28533, 28591, 32254, 29851, 
    28475, 29838, 25778, 24128, 19080, 15824, 12627, 9905, 5344, 1209, -5202, 
    -8103, -12054, -15205, -20255, -23137, -26681, -28947, -30337, -29454, 
    -30478, -30206, -30147, -29549, -25833, -23619, -20294, -17790, -13956, 
    -8757, -6131, -519, 3586, 6797, 11620, 15356, 19852, 21880, 25066, 28011, 
    29035, 30687, 30294, 30323, 28550, 28507, 26053, 23798, 20002, 18183, 
    14987, 9734, 4842, 1517, -2385, -7435, -11667, -15139, -19499, -21972, 
    -25424, -28032, -28110, -31344, -31331, -30018, -30865, -29366, -27092, 
    -24054, -20671, -16582, -12808, -9056, -6301, -2416, 4083, 7489, 11072, 
    16421, 19774, 22491, 24594, 27078, 29455, 30552, 31422, 29545, 29875, 
    28264, 26078, 25809, 22758, 19236, 13863, 9600, 5158, 177, -2435, -6452, 
    -10549, -13574, -17760, -21289, -24437, -25800, -28657, -30012, -30856, 
    -31555, -29812, -28218, -25638, -24357, -22126, -18032, -14958, -10740, 
    -6738, -2011, 3526, 6755, 11670, 13641, 19057, 21628, 23738, 27623, 
    28892, 30822, 31450, 32199, 29711, 27845, 28375, 24244, 21521, 18028, 
    13580, 11033, 6307, 1234, -1704, -6784, -10902, -15723, -19889, -22393, 
    -25997, -27172, -27386, -30259, -30722, -31350, -31470, -28013, -27197, 
    -25473, -21244, -20101, -14925, -12044, -7850, -3446, 1312, 6951, 11565, 
    14252, 19464, 20619, 24033, 27446, 28765, 28713, 30883, 31595, 30780, 
    29423, 28468, 24996, 22458, 17637, 14844, 9266, 6928, 1204, -3087, -5806, 
    -8787, -15275, -17372, -22005, -23097, -26408, -29684, -30489, -30380, 
    -30234, -31363, -28765, -27271, -26709, -22198, -18028, -14752, -9949, 
    -5494, -3910, 2173, 6940, 9565, 14831, 17151, 21780, 23278, 26676, 28989, 
    28371, 31312, 30024, 30162, 28110, 27346, 23852, 21461, 19032, 16039, 
    10664, 7758, 2876, -646, -5932, -9605, -13138, -17168, -21031, -26101, 
    -27311, -28736, -29069, -31836, -29730, -30319, -28648, -29030, -25531, 
    -21359, -19428, -16161, -11147, -6205, -2411, 1182, 7153, 9819, 12413, 
    17304, 22293, 22647, 27703, 27573, 29398, 29455, 29479, 29085, 28190, 
    27887, 24916, 22206, 18384, 15970, 10828, 6857, 3364, 298, -4931, -9055, 
    -15307, -18557, -20255, -23785, -27010, -28514, -29224, -31321, -30892, 
    -29768, -30344, -26738, -25630, -23493, -19082, -15121, -12422, -7928, 
    -3234, -606, 4443, 8531, 13198, 17226, 19275, 23629, 26889, 27499, 28514, 
    32017, 31616, 30574, 29712, 28871, 25499, 22616, 19389, 16130, 12997, 
    7928, 3042, -467, -4240, -9594, -13723, -17681, -20372, -22629, -25466, 
    -28422, -28892, -30885, -31675, -31441, -28468, -26551, -26037, -23470, 
    -20836, -16367, -12579, -8435, -2387, 1474, 5872, 9343, 13564, 18063, 
    20160, 24433, 25203, 29501, 28502, 29317, 31389, 30779, 30153, 28212, 
    25784, 24174, 19872, 16638, 12956, 8755, 4293, -1630, -6095, -8202, 
    -12296, -16454, -20581, -22436, -25772, -27807, -28535, -31012, -32568, 
    -29748, -30503, -28961, -26262, -23438, -21138, -17270, -13241, -8425, 
    -3661, 1214, 5121, 7136, 13604, 16624, 19587, 23733, 24774, 26320, 29163, 
    28619, 29639, 31206, 29449, 27646, 26368, 23250, 19268, 15593, 12580, 
    8544, 3928, 1426, -5308, -9924, -12632, -16404, -19603, -23557, -25197, 
    -29064, -27788, -29592, -29110, -29924, -31575, -27251, -26107, -23264, 
    -20249, -17500, -12324, -9247, -6068, -427, 3087, 8266, 12738, 16148, 
    20488, 23878, 24969, 27558, 29471, 30665, 31583, 31008, 30715, 27219, 
    25284, 23325, 19790, 15709, 13486, 8989, 4566, 441, -4867, -8826, -11883, 
    -14974, -19122, -22917, -26179, -27588, -30359, -31070, -30154, -29743, 
    -30534, -29781, -25946, -25087, -20356, -17467, -13545, -9187, -5323, 
    -1077, 2720, 9501, 10609, 17143, 19706, 22003, 25733, 27682, 29223, 
    30954, 31230, 30466, 30691, 29013, 26226, 23408, 21287, 18803, 14067, 
    8988, 6069, 2255, -2864, -8350, -10821, -15871, -19953, -22210, -26393, 
    -27489, -29989, -30812, -31913, -30850, -29039, -30269, -27506, -24726, 
    -20253, -17302, -13140, -9949, -5558, -1236, 3417, 7586, 11430, 15525, 
    18396, 21987, 24644, 27965, 30199, 30262, 30280, 30100, 31137, 28714, 
    24890, 25398, 21434, 17852, 13812, 10565, 6242, 10, -1282, -7127, -10707, 
    -14675, -18676, -22945, -24890, -26704, -29926, -29140, -29440, -31153, 
    -29157, -29092, -27350, -23031, -20274, -18210, -14202, -10023, -6257, 
    -1294, 2656, 8292, 12274, 15808, 18345, 22646, 25110, 28794, 29081, 
    29140, 29335, 29272, 28331, 28078, 25950, 23467, 23227, 17712, 15214, 
    10673, 6851, 2111, -1673, -6681, -10684, -14049, -18379, -22025, -24795, 
    -25904, -27920, -30267, -30503, -29374, -29534, -27866, -26391, -24104, 
    -21827, -18533, -14369, -10189, -5204, -972, 1060, 5846, 10306, 14656, 
    17774, 20947, 24684, 27302, 29313, 29684, 30282, 30167, 29301, 29423, 
    26466, 24067, 22538, 18454, 15458, 10021, 7511, 2431, -3251, -6016, 
    -9506, -14207, -18491, -23306, -24861, -26233, -28884, -30080, -31102, 
    -30066, -29806, -28400, -28255, -26232, -23566, -19971, -15327, -9808, 
    -5825, -1181, 3083, 4633, 9559, 15065, 16422, 22543, 24228, 26214, 29147, 
    29053, 30412, 31538, 30648, 29624, 28017, 24613, 20465, 19537, 15132, 
    9745, 6848, 4441, -1492, -4451, -9731, -13550, -16789, -20532, -25102, 
    -27531, -26979, -29668, -30338, -31632, -29681, -30191, -26426, -24973, 
    -21919, -18769, -15329, -11351, -7506, -4435, 1654, 5424, 9693, 12817, 
    18155, 20710, 24963, 26612, 26696, 28046, 29675, 29762, 29915, 29188, 
    26913, 24749, 23528, 17729, 14760, 11497, 7073, 4032, -805, -4934, 
    -10701, -13710, -17676, -19603, -23191, -27044, -28976, -29908, -30203, 
    -30384, -30427, -30344, -26907, -24495, -23768, -18762, -15801, -11830, 
    -8092, -4089, 1210, 4719, 9849, 13568, 17563, 21452, 25031, 26074, 28398, 
    29482, 29643, 29116, 30640, 29164, 27282, 25443, 22005, 20036, 16722, 
    11182, 8355, 4893, -483, -4269, -9822, -13383, -17681, -20520, -23011, 
    -26391, -29514, -28461, -30052, -30913, -29108, -27876, -26630, -26086, 
    -24626, -19632, -16771, -12185, -8758, -5162, -560, 5271, 10058, 12523, 
    17160, 19506, 23314, 26044, 27830, 28309, 30085, 32136, 31388, 29519, 
    28381, 25659, 24130, 19252, 16935, 11695, 8514, 4261, -591, -5169, -8185, 
    -14341, -16653, -21201, -22305, -27367, -27674, -30881, -29311, -31673, 
    -30762, -30437, -27359, -24914, -22292, -19261, -16667, -11633, -9703, 
    -4800, -387, 2799, 8279, 12476, 16899, 18606, 24757, 27041, 28745, 28451, 
    30852, 31436, 29828, 28975, 26996, 24391, 23752, 21488, 15499, 13734, 
    8102, 5382, 1393, -3561, -8911, -12355, -17823, -19831, -24147, -26267, 
    -26537, -29161, -30686, -30504, -31925, -30423, -26737, -26721, -23206, 
    -20471, -16507, -12206, -8250, -6329, 1074, 3322, 6670, 14186, 16796, 
    20128, 21841, 25344, 26803, 29995, 31347, 30181, 30217, 30186, 27092, 
    26068, 23843, 20733, 17144, 13956, 9121, 6174, 1808, -3558, -8216, 
    -11946, -14723, -19649, -21684, -24266, -29347, -29344, -30246, -30622, 
    -31866, -30175, -27329, -26117, -24044, -20721, -18706, -14044, -9092, 
    -4561, -1057, 3049, 7658, 12063, 15182, 19035, 22242, 26661, 27752, 
    29528, 31453, 29057, 30969, 28871, 27641, 26061, 22608, 21525, 17566, 
    14279, 9403, 4880, 933, -3794, -8327, -10521, -15531, -18660, -22218, 
    -24663, -28368, -29105, -31314, -31554, -30675, -28781, -28642, -26193, 
    -24867, -19827, -18642, -15097, -9758, -6651, -1102, 2817, 7575, 10772, 
    14243, 18777, 21576, 26290, 28178, 29675, 30032, 30228, 29229, 31644, 
    27425, 24844, 24377, 22268, 16522, 15150, 10092, 5259, 1016, -3655, 
    -7563, -10187, -15420, -19287, -23220, -24793, -27292, -28843, -31645, 
    -30276, -29798, -30738, -29365, -25559, -25291, -20361, -18054, -15169, 
    -9897, -6725, -1586, 2558, 7301, 12195, 15367, 18494, 22298, 23772, 
    26891, 28723, 30704, 31091, 30774, 28621, 29363, 26137, 24730, 21379, 
    18729, 14166, 10978, 5718, 1863, -4176, -6461, -10648, -14089, -19057, 
    -21837, -25916, -27191, -29670, -30503, -30622, -31117, -29850, -28141, 
    -27259, -25011, -20775, -17548, -14624, -11319, -5737, -3304, 1135, 6874, 
    9665, 15930, 17208, 21030, 25396, 28028, 29222, 31605, 29219, 30307, 
    29702, 28807, 26765, 26255, 21005, 18782, 13925, 11190, 7411, 1745, 
    -1646, -6604, -10329, -16304, -19270, -21010, -26084, -26565, -27982, 
    -30423, -31772, -30671, -30539, -28709, -26801, -24821, -22608, -17387, 
    -15534, -10753, -6540, -1755, 1534, 7389, 10886, 13390, 17560, 20649, 
    24835, 26199, 28558, 30194, 30695, 30104, 30389, 30502, 27438, 24639, 
    22486, 18577, 15787, 11327, 6299, 1741, -1147, -6052, -9954, -15415, 
    -18617, -22489, -25179, -27690, -29967, -29711, -30872, -30365, -30738, 
    -29999, -27854, -26180, -22650, -18740, -15519, -10584, -7482, -3426, 
    1927, 6582, 9825, 14706, 17373, 22489, 24117, 26103, 28531, 29527, 30746, 
    30986, 29602, 30075, 27468, 25398, 21337, 19028, 15088, 11230, 6096, 
    3749, -1404, -4974, -8819, -12356, -16971, -20301, -24582, -26002, 
    -27713, -31001, -31915, -30733, -30587, -30295, -27370, -25413, -23059, 
    -19604, -15696, -12582, -6223, -3759, 1848, 5580, 10601, 14194, 16292, 
    19964, 23023, 26710, 28848, 30440, 28885, 30569, 29502, 28087, 28737, 
    25129, 23096, 20975, 15309, 13098, 7419, 4107, -1516, -5934, -9340, 
    -11807, -17765, -21942, -25411, -27112, -28293, -28912, -29912, -31948, 
    -29913, -29967, -28375, -23974, -22537, -20914, -17448, -12111, -7923, 
    -4436, 64, 5459, 8117, 13645, 18038, 20871, 23512, 24358, 27946, 29068, 
    29969, 30760, 30961, 29974, 27521, 27235, 23736, 19803, 16488, 12451, 
    8106, 4257, -400, -4955, -10404, -12999, -15266, -19511, -23328, -27452, 
    -26956, -31221, -30461, -31438, -32049, -30778, -27992, -25567, -23547, 
    -21501, -17715, -12270, -8634, -3939, -243, 3316, 9033, 12793, 16644, 
    20630, 22047, 25106, 27186, 29434, 29192, 29192, 30474, 28037, 29134, 
    26111, 22621, 20942, 16753, 11927, 8869, 5346, 1347, -4435, -9014, 
    -12676, -17336, -19637, -23292, -26442, -29418, -30008, -30984, -29775, 
    -30631, -29851, -27322, -25996, -24462, -21283, -16474, -13259, -10301, 
    -4181, -390, 3387, 9497, 12932, 15246, 19726, 22773, 25497, 26800, 30287, 
    29672, 31585, 30201, 29573, 29050, 25791, 23293, 19904, 17265, 13226, 
    8774, 4291, 1053, -5167, -8205, -10493, -14271, -19473, -23696, -25580, 
    -27958, -27687, -31575, -31184, -29934, -29695, -28214, -26802, -23871, 
    -21073, -16884, -13854, -9014, -5904, -1981, 2434, 7358, 10290, 15198, 
    19290, 23026, 23924, 27192, 28950, 30366, 32491, 31958, 30101, 28539, 
    25089, 24088, 20694, 16935, 14394, 9910, 4913, 814, -4705, -8006, -11002, 
    -16126, -20098, -22348, -24101, -28560, -28557, -30801, -30975, -30709, 
    -31188, -28571, -26095, -23398, -20923, -18174, -15376, -9029, -6561, 
    -1247, 1842, 6135, 12280, 16427, 20080, 21661, 25691, 25845, 30488, 
    31017, 30573, 30748, 28874, 28417, 25563, 23797, 20703, 16406, 14384, 
    9956, 7199, 2256, -3953, -8501, -12514, -16697, -19043, -22975, -24863, 
    -28010, -28883, -29748, -30642, -30100, -30948, -29807, -27330, -23270, 
    -22846, -16787, -14418, -12001, -6430, -1364, 3691, 6834, 10484, 15295, 
    17101, 23029, 24263, 27359, 29213, 30762, 29754, 31104, 30281, 30103, 
    27358, 22953, 22336, 17617, 13262, 11711, 5802, 2710, -2599, -7576, 
    -12015, -14318, -18833, -22739, -25160, -26436, -28844, -30735, -30139, 
    -29833, -30873, -29237, -27212, -24180, -20407, -17712, -15540, -10587, 
    -5492, -1917, 2446, 7046, 11440, 15616, 18976, 21001, 24778, 27739, 
    28560, 30152, 30203, 31865, 29235, 28397, 28402, 24641, 22744, 19051, 
    15801, 12745, 5541, 2580, -860, -4973, -10551, -13751, -18523, -21647, 
    -23562, -26764, -29422, -28737, -32291, -31277, -30634, -28508, -27408, 
    -25750, -21852, -19112, -15276, -11701, -6647, -2495, 1436, 7349, 10637, 
    13920, 18286, 21404, 24331, 25401, 29376, 28812, 30462, 29890, 29099, 
    29049, 27065, 25086, 22538, 18211, 15161, 10061, 7265, 2503, 228, -6831, 
    -11328, -12974, -17403, -20772, -25317, -26845, -29781, -30493, -32164, 
    -31003, -30404, -28903, -27287, -25493, -21249, -20741, -15783, -11647, 
    -7737, -2826, 1625, 5538, 10659, 13362, 17732, 21203, 24802, 27812, 
    27438, 30352, 29101, 31071, 31921, 28924, 28162, 25167, 22341, 19493, 
    14947, 12114, 6841, 1971, -1962, -5438, -8586, -13803, -17213, -20961, 
    -22951, -25721, -27056, -31362, -32150, -30413, -30170, -29081, -28846, 
    -24065, -22575, -21208, -15656, -12580, -7668, -3452, -366, 4010, 9739, 
    13851, 17002, 20242, 23818, 26535, 28002, 29351, 29780, 31706, 30136, 
    28695, 27127, 25863, 22732, 20158, 17755, 11396, 7243, 3283, -1255, 
    -4186, -9995, -13557, -17104, -20087, -24016, -26446, -28318, -29576, 
    -30380, -32275, -29545, -29129, -28481, -25207, -21545, -19587, -14833, 
    -12205, -7173, -4919, -1141, 4961, 9238, 13337, 16591, 18884, 24674, 
    26221, 28733, 28903, 32217, 30468, 30805, 29533, 28673, 27116, 23728, 
    19154, 17094, 11024, 8807, 5315, -1901, -4136, -7056, -14698, -16826, 
    -20502, -24890, -25816, -28012, -31257, -30949, -29952, -29985, -31225, 
    -26759, -26426, -22913, -21432, -16098, -13437, -10089, -3562, -1251, 
    3185, 8984, 12491, 17272, 21002, 22437, 26459, 29392, 28555, 30432, 
    30193, 30801, 29286, 28047, 26212, 21816, 19634, 18002, 11914, 8679, 
    4566, 564, -4661, -8197, -13571, -16538, -19493, -22007, -25951, -26723, 
    -30682, -31340, -30166, -29745, -29092, -28936, -25727, -25199, -19978, 
    -17353, -13139, -9544, -5293, -879, 3647, 7960, 11157, 15212, 19001, 
    22601, 24535, 27403, 31186, 29956, 31389, 30354, 29846, 28702, 25384, 
    22052, 19298, 16352, 13117, 9536, 5434, 1064, -4588, -8195, -12975, 
    -17099, -19652, -23558, -26934, -27082, -29865, -29761, -31536, -30962, 
    -31028, -28495, -26876, -23418, -20614, -17973, -12740, -9629, -4863, 
    -1822, 3560, 8379, 12055, 15979, 21091, 22348, 25453, 28512, 29964, 
    31515, 31099, 30589, 30422, 28416, 27275, 24419, 19711, 18472, 13598, 
    10288, 4751, 1193, -3827, -6699, -11882, -15008, -18339, -22816, -23806, 
    -26277, -29503, -31003, -30828, -29752, -30910, -30031, -27672, -23941, 
    -21120, -17891, -13789, -8675, -4491, -2194, 3172, 7629, 12361, 15100, 
    19790, 22395, 26233, 25839, 27854, 29755, 30996, 30562, 30048, 28239, 
    26012, 23291, 21513, 17550, 13509, 9938, 6902, 1657, -3539, -7777, 
    -11175, -15328, -19043, -22473, -25464, -28502, -28177, -29509, -31617, 
    -32028, -30215, -27907, -28121, -24862, -19616, -17157, -13983, -10242, 
    -5782, -1330, 2433, 7218, 12292, 14997, 18239, 20883, 24969, 28983, 
    29434, 30940, 31385, 31574, 29601, 29274, 26985, 23903, 21101, 18112, 
    15006, 8981, 5466, 1978, -2892, -6367, -10193, -15931, -17938, -20596, 
    -25411, -26770, -29788, -31745, -30124, -30969, -29461, -28166, -27450, 
    -26002, -21040, -17910, -13415, -11246, -6000, -1285, 3008, 7619, 9579, 
    14262, 19088, 22311, 25523, 26570, 30288, 29345, 30548, 31320, 29441, 
    29003, 27219, 23366, 20423, 17281, 14792, 10343, 7077, 3607, -211, -6291, 
    -9555, -15579, -18134, -22332, -23553, -26048, -28197, -30502, -30690, 
    -31594, -29814, -28173, -27435, -23859, -20797, -19104, -15467, -11976, 
    -6491, -3003, 106, 4582, 10975, 15869, 16823, 22679, 24239, 27999, 29220, 
    29795, 29438, 31110, 30474, 28765, 26403, 24217, 22670, 18567, 15616, 
    12028, 6247, 2834, -2366, -5734, -10609, -14681, -19167, -21010, -23209, 
    -26037, -29243, -30206, -30637, -31134, -31322, -27839, -28429, -26468, 
    -21935, -19445, -14589, -12975, -6060, -2950, 1008, 6345, 10214, 13521, 
    18702, 21343, 23378, 26936, 30278, 30861, 31996, 30973, 30811, 29093, 
    27679, 24172, 23617, 19929, 15890, 10977, 6325, 4590, 312, -6511, -9513, 
    -14614, -18606, -20531, -22773, -25855, -28567, -29969, -28930, -30970, 
    -29674, -27712, -27837, -25996, -23642, -18919, -15655, -12421, -8414, 
    -3855, 370, 5644, 8262, 12503, 16686, 20734, 22699, 26553, 28740, 28949, 
    31376, 32038, 29738, 30405, 28253, 26779, 21900, 20769, 14391, 10304, 
    8891, 4671, -1587, -4403, -9322, -13649, -18076, -21322, -23412, -27225, 
    -28780, -28476, -29518, -31597, -30952, -29521, -26844, -24295, -23853, 
    -18809, -16886, -13693, -8729, -2611, 1672, 3715, 9733, 13113, 17120, 
    21680, 24136, 27328, 27713, 29660, 30686, 30669, 31192, 29305, 26995, 
    26291, 22974, 18730, 16409, 12456, 8491, 4500, -778, -5235, -9204, 
    -13056, -16108, -20391, -23643, -26510, -27966, -29383, -29583, -29977, 
    -29927, -29415, -27899, -25899, -24270, -20308, -16571, -12063, -7906, 
    -5858, 1268, 2723, 7192, 11100, 17510, 20221, 22416, 26022, 28963, 29537, 
    30165, 31522, 29267, 29958, 29627, 25137, 23164, 19606, 16083, 13801, 
    8242, 4048, -174, -4511, -7785, -13998, -15130, -19622, -24123, -26663, 
    -28123, -27764, -29674, -31019, -31604, -29175, -26873, -25696, -24210, 
    -19691, -16399, -14905, -7888, -5265, 1082, 3535, 7693, 13178, 17772, 
    21397, 24318, 25851, 27177, 28400, 31408, 30988, 30139, 29720, 28139, 
    25592, 22359, 19574, 17133, 14325, 9730, 3973, 577, -4466, -6939, -12962, 
    -15309, -20964, -23195, -26336, -28511, -30068, -28769, -30364, -30501, 
    -30439, -27070, -26193, -24667, -21490, -17487, -13794, -9383, -3796, 
    -536, 2986, 8335, 13150, 15426, 19531, 22754, 24765, 28986, 29558, 31358, 
    31235, 30779, 29526, 28316, 24891, 22650, 21894, 16172, 15144, 10151, 
    5323, 524, -4397, -6391, -11276, -16658, -18225, -22638, -25026, -27287, 
    -29872, -29547, -32658, -29274, -31351, -28470, -26177, -23129, -21030, 
    -16908, -13478, -10099, -5564, -2908, 4298, 8228, 12294, 13967, 18832, 
    20897, 26587, 26789, 29778, 29435, 30451, 30198, 30208, 28207, 27317, 
    22563, 22058, 18570, 15547, 8715, 6832, 2110, -1195, -6535, -11511, 
    -13873, -18483, -22265, -24835, -27500, -28827, -30537, -31425, -30630, 
    -29503, -29099, -27293, -24433, -20537, -16366, -12713, -9278, -6153, 
    -1493, 3659, 6395, 12019, 15139, 18532, 22790, 26389, 26542, 28250, 
    30273, 32024, 30490, 30262, 29115, 26678, 24420, 21587, 18854, 15374, 
    10599, 5588, 1783, -2021, -5942, -10482, -14943, -19310, -22734, -24911, 
    -26078, -28922, -30414, -30264, -31659, -29288, -28843, -25598, -24903, 
    -22348, -17738, -14763, -10782, -6757, -2390, 1600, 6935, 11868, 14649, 
    18910, 21499, 24535, 26439, 27262, 30450, 29920, 29632, 28956, 28640, 
    27136, 23734, 21915, 17543, 14980, 11000, 6961, 1487, -2484, -7108, 
    -10226, -15582, -19485, -23066, -24175, -26640, -29128, -30840, -29516, 
    -30321, -30277, -29867, -26915, -24171, -20723, -19117, -15064, -11110, 
    -7421, -2339, 285, 6237, 10943, 14881, 17123, 21804, 24690, 28186, 30459, 
    29965, 30508, 31257, 30911, 28763, 26664, 25315, 21662, 20016, 16643, 
    11719, 8758, 2173, -2240, -5209, -10034, -14933, -18583, -20561, -24521, 
    -27499, -28364, -30068, -28994, -30464, -29688, -27783, -27677, -25842, 
    -23257, -19104, -14611, -11226, -6604, -2249, 2237, 4953, 8823, 13785, 
    16135, 21557, 25520, 26357, 28937, 29653, 31131, 30668, 30736, 29857, 
    27182, 23914, 21216, 19337, 15767, 12020, 6282, 4608, -1634, -6480, 
    -8673, -12343, -16997, -20924, -22847, -25732, -26998, -28703, -31175, 
    -31800, -31189, -28582, -27371, -25015, -24207, -19654, -16382, -11387, 
    -8996, -3722, 828, 5890, 7952, 14673, 17645, 19775, 25506, 26473, 29636, 
    30045, 31229, 31403, 30246, 30032, 26751, 25185, 22924, 19405, 14934, 
    12573, 8568, 3867, -779, -6282, -9058, -14327, -18423, -19725, -23004, 
    -25598, -28839, -30104, -31300, -30059, -28898, -29126, -27850, -25458, 
    -22992, -19677, -16379, -12274, -8558, -4126, 1365, 5579, 7762, 12221, 
    18387, 20362, 23371, 25630, 26866, 29739, 31340, 30276, 29896, 29821, 
    28753, 25361, 23028, 18757, 16082, 13123, 7473, 4705, 895, -4571, -9788, 
    -12871, -17269, -19337, -22967, -26074, -28049, -29626, -29309, -31256, 
    -28819, -31166, -27306, -26183, -23768, -20797, -16555, -12733, -8973, 
    -3788, -1061, 4798, 9970, 12919, 15667, 21740, 23888, 25697, 29707, 
    31064, 29634, 31039, 29486, 28617, 27278, 25413, 24502, 19150, 16088, 
    13521, 8495, 3415, 703, -4367, -8842, -12806, -15710, -21075, -23863, 
    -24429, -29619, -29606, -30628, -29508, -29926, -28617, -28334, -25971, 
    -23797, -19988, -16846, -13830, -7659, -3997, 483, 3077, 7844, 12347, 
    16324, 19593, 21776, 26593, 28686, 29711, 29653, 30372, 30280, 30338, 
    28929, 25311, 24125, 21987, 17408, 14287, 8612, 6135, -54, -4868, -7743, 
    -13036, -15954, -19783, -22011, -26093, -27533, -29558, -29927, -30026, 
    -31024, -28393, -28986, -26458, -23708, -22127, -17391, -13675, -9426, 
    -5454, -2237, 4322, 8027, 10773, 14067, 20796, 22080, 24895, 26106, 
    31096, 30063, 30599, 30849, 29162, 27520, 25535, 24335, 20379, 18803, 
    14756, 8635, 5832, 948, -4785, -6518, -11549, -14952, -18331, -22801, 
    -25892, -28140, -28543, -30363, -31804, -30295, -30891, -29866, -25992, 
    -24616, -19999, -17378, -14386, -9500, -7226, -1810, 4548, 7159, 10809, 
    14964, 19918, 21164, 25587, 26998, 29279, 29455, 30520, 30168, 29774, 
    28811, 28136, 23241, 21809, 17240, 14596, 11452, 5459, 1671, -2261, 
    -6888, -10939, -15126, -19279, -22048, -24726, -27368, -27999, -30262, 
    -30207, -31183, -28451, -28097, -27568, -23808, -21439, -18242, -13999, 
    -10103, -4257, -1233, 2368, 6907, 12633, 15747, 19959, 22223, 26097, 
    27665, 30131, 30684, 31327, 30256, 30196, 30052, 27583, 25485, 21744, 
    17066, 14866, 10084, 5647, 3444, -3059, -6246, -10797, -14210, -18976, 
    -22788, -25367, -27278, -29235, -29730, -29772, -31265, -29580, -29274, 
    -27819, -24491, -22511, -17628, -14409, -10290, -4761, -3488, 1269, 5157, 
    10650, 14724, 17596, 23083, 25117, 27051, 29311, 31105, 30366, 30535, 
    29377, 30140, 26379, 23515, 21420, 17347, 14683, 12176, 7450, 2652, 
    -2016, -7664, -10302, -15015, -19619, -21482, -22900, -27867, -29471, 
    -29963, -30288, -31033, -31182, -28801, -27880, -24675, -22030, -17468, 
    -16195, -11823, -7324, -3599, 1671, 6190, 9134, 14393, 19055, 21019, 
    25107, 27921, 28602, 29812, 29944, 31431, 30453, 27632, 26882, 24966, 
    21865, 18122, 17132, 9582, 6829, 3327, -1919, -7059, -9373, -14301, 
    -18504, -21910, -22886, -27094, -28082, -31101, -30849, -29582, -30135, 
    -28706, -27226, -25960, -22939, -18915, -13921, -9987, -7627, -2499, 268, 
    7015, 10140, 15810, 18564, 20962, 24604, 27810, 28466, 30506, 30133, 
    31652, 31812, 29933, 28463, 25186, 21297, 18430, 15253, 11604, 6152, 
    2041, 170, -4173, -10274, -13511, -17168, -22337, -23041, -27257, -27482, 
    -30588, -30502, -30467, -29541, -29654, -25797, -27264, -22505, -19724, 
    -15261, -12103, -7603, -1990, 2500, 6570, 10674, 14410, 17138, 21867, 
    23640, 25060, 27877, 30274, 30778, 30822, 31310, 28954, 28070, 23941, 
    23698, 19648, 16414, 11665, 9657, 3407, -1091, -4322, -8083, -14444, 
    -17434, -20663, -22655, -26284, -28693, -29769, -31339, -32536, -29898, 
    -29313, -28526, -24865, -22456, -17929, -15899, -11807, -9525, -4056, 
    1488, 4695, 9087, 14800, 17548, 21985, 22834, 26312, 27545, 31221, 31094, 
    29676, 31931, 28760, 28073, 26094, 23588, 20601, 15651, 13743, 8700, 
    3997, -795, -3129, -8821, -13471, -17925, -20055, -24691, -27019, -29305, 
    -29312, -30391, -30929, -30490, -28944, -27053, -26545, -24049, -19920, 
    -17656, -12438, -8646, -4829, 1197, 4518, 9028, 13914, 16869, 21758, 
    22035, 26277, 26855, 30189, 30711, 31711, 31424, 29980, 28091, 26266, 
    23353, 21888, 17135, 11669, 9282, 4935, 1232, -4800, -9226, -13720, 
    -14977, -21460, -22837, -25596, -27791, -29026, -29527, -30265, -31240, 
    -28830, -28545, -25398, -23607, -21777, -18005, -13956, -7704, -4606, 
    223, 2696, 9327, 12913, 16037, 20355, 24256, 23990, 28042, 29433, 30234, 
    30758, 30867, 29274, 27970, 26035, 22868, 19995, 18206, 12656, 10518, 
    4558, 520, -3934, -8083, -12499, -17603, -18556, -22084, -25582, -26334, 
    -30078, -30261, -31057, -31192, -28090, -28668, -26586, -22179, -20240, 
    -17485, -13946, -8579, -4726, -1559, 4421, 8925, 12975, 15291, 19525, 
    21688, 26879, 28283, 29269, 31324, 31089, 31115, 29976, 28350, 27328, 
    24193, 20378, 18206, 13686, 9797, 6151, 1125, -2836, -8341, -10573, 
    -16341, -18437, -22853, -25383, -28328, -29954, -29077, -30263, -29396, 
    -28848, -27781, -26025, -23994, -20297, -17951, -14983, -10274, -4947, 
    -747, 4928, 7435, 10660, 14997, 19169, 23931, 25218, 26794, 29977, 30451, 
    30130, 30685, 30874, 28805, 27271, 24120, 20897, 17085, 14339, 11374, 
    5746, 1143, -4019, -8047, -12196, -14747, -18099, -23106, -25592, -28586, 
    -27586, -28755, -32008, -30182, -31171, -30134, -26449, -23753, -21865, 
    -17390, -12983, -11273, -7141, -2221, 3522, 7166, 12180, 15956, 20218, 
    23594, 24390, 25645, 29323, 29666, 29841, 30917, 30052, 29360, 26170, 
    25657, 20025, 19362, 13583, 11129, 4712, 1048, -3207, -7316, -10109, 
    -14745, -18333, -22890, -25126, -25404, -28998, -30780, -29665, -31423, 
    -30453, -27996, -26769, -25508, -20557, -18824, -15244, -10436, -7798, 
    -2320, 1600, 6876, 10281, 13409, 17293, 21620, 24189, 26188, 27377, 
    31326, 30096, 30980, 30187, 27674, 27211, 23789, 20698, 18188, 15815, 
    11965, 8260, 3758, -2258, -6068, -11816, -14133, -16725, -21581, -25670, 
    -27295, -30105, -30146, -31152, -30772, -30817, -29036, -27475, -25089, 
    -22555, -18352, -16200, -12261, -8524, -1640, 178, 4766, 9220, 13881, 
    18100, 21057, 24855, 26954, 28895, 30402, 31322, 30104, 29760, 29294, 
    25988, 23747, 21997, 19683, 15015, 11472, 7893, 2576, -3131, -6136, 
    -9998, -14259, -18637, -21468, -24897, -25208, -27195, -30116, -30327, 
    -30450, -29853, -29768, -26777, -24125, -23032, -18893, -14459, -11268, 
    -7589, -2762, 2745, 6817, 10386, 14596, 17626, 22264, 22891, 24933, 
    27725, 29611, 30800, 31316, 31270, 28314, 26706, 23865, 23976, 20214, 
    15351, 12466, 8090, 3607, -410, -4153, -9755, -14623, -17564, -22067, 
    -23811, -27449, -29857, -30235, -31306, -30846, -31056, -30285, -26980, 
    -25101, -21992, -19205, -14805, -11844, -7492, -4596, 2121, 5491, 9100, 
    13521, 18509, 19606, 23900, 26103, 29596, 28806, 30155, 31070, 31469, 
    30285, 26851, 25110, 22262, 20038, 16320, 11643, 7801, 4945, -1503, 
    -4338, -7771, -13762, -18757, -20794, -22913, -27040, -27745, -28439, 
    -30557, -30451, -29541, -30067, -27721, -26915, -23086, -18892, -15119, 
    -11638, -9426, -3043, -167, 4574, 8405, 13090, 17866, 20936, 23825, 
    26315, 27781, 29425, 30700, 31701, 30553, 29933, 28556, 24606, 21611, 
    19034, 16824, 13014, 8657, 4519, -702, -4591, -8872, -12572, -16671, 
    -21867, -22721, -25943, -29729, -29482, -30526, -30146, -29333, -30085, 
    -27481, -24800, -23233, -20036, -17109, -12671, -8222, -5711, -253, 4690, 
    9073, 13706, 16968, 20003, 22759, 24718, 26860, 28737, 30221, 32042, 
    31138, 29215, 28111, 26156, 23728, 19677, 16829, 11704, 9088, 5520, 1581, 
    -2472, -10043, -14240, -15653, -20439, -22843, -24779, -27751, -30537, 
    -30467, -30217, -30051, -29557, -29439, -26285, -24067, -19593, -16168, 
    -13484, -9155, -4419, -705, 3856, 8822, 12621, 14884, 18862, 22705, 
    25074, 29064, 29142, 30954, 31134, 28985, 29631, 28308, 26956, 24297, 
    21773, 16593, 12248, 9638, 3843, 489, -3639, -8240, -12986, -16152, 
    -18323, -23496, -24693, -27238, -28631, -31337, -31732, -31572, -30991, 
    -28429, -24876, -24459, -21699, -18892, -13424, -10254, -4493, -386, 
    3385, 6896, 12012, 17165, 18720, 22927, 24872, 27927, 29518, 29587, 
    29514, 30449, 29849, 26968, 27146, 25080, 22547, 17352, 13371, 9986, 
    4191, 1453, -3547, -6764, -12462, -14999, -20743, -23592, -25819, -27457, 
    -30548, -29532, -30642, -29463, -30139, -29426, -26709, -23231, -21322, 
    -18354, -15505, -10372, -5998, -313, 3600, 6193, 11047, 14926, 20018, 
    22563, 25390, 26684, 29652, 32016, 31973, 30571, 28723, 28329, 27208, 
    24168, 22040, 17614, 13633, 9400, 4607, 1478, -4628, -6546, -11569, 
    -15907, -19992, -21273, -26247, -25708, -30154, -28590, -31782, -30318, 
    -29771, -29624, -25205, -24309, -21439, -18453, -14158, -9950, -4867, 
    -2258, 2926, 7158, 11073, 15879, 20077, 20830, 25683, 27064, 30323, 
    28779, 30379, 31480, 29716, 28654, 26839, 23205, 22235, 18721, 14682, 
    10569, 5782, 2922, -900, -5718, -10223, -15171, -18433, -20763, -23383, 
    -27804, -28967, -30004, -32293, -30691, -28662, -28198, -26746, -24858, 
    -21530, -17906, -14615, -10340, -6196, -1983, 2341, 6998, 10568, 14663, 
    19969, 22565, 23877, 25357, 29006, 30227, 30714, 31200, 29337, 28584, 
    27200, 26384, 21782, 18238, 14272, 9366, 6272, 1561, -1949, -5486, -9759, 
    -15085, -17004, -20264, -25551, -26016, -30012, -30357, -30757, -31450, 
    -30516, -28775, -26309, -25290, -22128, -20031, -15814, -9719, -6908, 
    -2415, 1578, 6207, 11310, 15141, 19257, 21899, 23805, 25482, 28696, 
    31259, 31053, 31348, 30318, 29438, 26877, 25334, 21891, 18397, 14365, 
    11305, 8888, 1351, -1023, -6772, -9953, -14509, -17814, -21720, -25186, 
    -26074, -28268, -28644, -29091, -29341, -30027, -28798, -28273, -26156, 
    -22072, -17711, -15180, -13094, -8079, -3956, 641, 6807, 10424, 13346, 
    18005, 20436, 23665, 26312, 28747, 29974, 32074, 30795, 31012, 29051, 
    27038, 24340, 24003, 20489, 15126, 12563, 7167, 3461, 16, -5404, -10381, 
    -13534, -17506, -21628, -24995, -26094, -28814, -30224, -30983, -30380, 
    -30551, -30736, -26922, -25511, -24006, -19697, -15846, -13647, -8298, 
    -3088, 861, 6244, 9453, 14935, 16379, 19680, 23629, 25998, 26892, 30307, 
    31554, 30467, 31783, 30709, 26432, 26212, 23041, 18716, 16217, 11582, 
    8295, 4519, 246, -5275, -10363, -12796, -16662, -21777, -23797, -27053, 
    -28536, -29841, -31155, -30711, -29207, -30478, -28221, -24554, -22901, 
    -19052, -14915, -13420, -7229, -5047, -371, 4372, 7388, 13279, 17628, 
    20737, 23237, 25818, 28554, 28618, 31979, 29906, 31187, 30227, 29458, 
    25424, 23532, 18879, 17600, 12442, 8870, 4098, 974, -4794, -7418, -13276, 
    -18020, -21031, -24212, -26287, -27454, -30143, -30328, -30994, -29671, 
    -29526, -27401, -25971, -22246, -20424, -17461, -11465, -7732, -3939, 
    -1758, 4148, 8758, 13696, 16992, 21600, 22216, 25742, 28460, 30890, 
    30166, 29161, 29463, 29755, 28526, 26066, 24136, 21550, 15969, 12159, 
    9084, 3946, 708, -5181, -9833, -12706, -17412, -19263, -23362, -27003, 
    -28915, -27637, -29330, -29876, -32149, -30168, -27816, -26936, -23526, 
    -19184, -18016, -11909, -8732, -4179, -449, 4054, 7917, 12538, 15380, 
    19783, 22731, 25381, 26736, 30586, 29729, 32150, 31510, 29712, 28656, 
    26235, 23056, 22281, 16254, 12804, 8904, 4781, 1320, -3712, -6928, 
    -12169, -14621, -19827, -21536, -24971, -26618, -30220, -31437, -31578, 
    -29651, -31165, -27285, -26195, -23965, -21885, -17467, -13050, -8310, 
    -5457, -712, 3628, 7824, 12671, 17012, 18339, 23394, 26355, 27064, 28763, 
    29743, 32026, 29968, 29957, 28854, 27226, 24926, 21026, 17341, 13682, 
    9610, 6486, 83, -3002, -7875, -11541, -15004, -18922, -23571, -24835, 
    -29084, -28565, -29676, -30631, -31967, -29742, -28198, -25827, -24460, 
    -20557, -17177, -14473, -9213, -5715, -1703, 2708, 7249, 11291, 14931, 
    17802, 22495, 26422, 28481, 28433, 30407, 31073, 30557, 30473, 28265, 
    26677, 23882, 21367, 16791, 12738, 9013, 5877, 2636, -3276, -7104, 
    -11219, -14111, -18742, -23236, -25843, -26299, -28230, -29577, -30146, 
    -31822, -29874, -28704, -27627, -24413, -19963, -17439, -14890, -11236, 
    -6526, -1284, 4038, 6916, 10574, 14866, 17362, 20750, 24771, 28370, 
    28449, 30439, 28977, 30279, 29619, 27934, 26804, 25006, 21487, 18908, 
    13312, 9775, 5648, 2414, -2892, -6591, -10478, -13890, -19765, -21120, 
    -23570, -26807, -27839, -29671, -31406, -31768, -29723, -27990, -28063, 
    -24802, -22573, -18370, -14375, -9948, -7313, -2263, 1822, 7393, 12277, 
    15900, 17476, 21623, 24905, 26918, 30511, 29832, 32034, 30142, 29670, 
    28235, 28496, 24496, 22134, 17101, 16816, 11744, 7282, 2327, -1310, 
    -5570, -10182, -14101, -19325, -21651, -23831, -27264, -28843, -29660, 
    -29789, -30746, -30899, -30066, -27310, -25923, -21814, -19361, -15148, 
    -11426, -5886, -3568, 866, 4557, 11862, 13924, 18141, 21436, 23410, 
    27184, 28179, 30175, 30732, 29881, 30221, 29649, 26925, 26241, 22451, 
    18480, 14903, 11507, 7358, 2959, -592, -4353, -10172, -13946, -16531, 
    -20873, -24014, -27180, -28296, -29382, -30607, -30568, -30736, -30598, 
    -27099, -25623, -23015, -18982, -15049, -12498, -9162, -3580, 244, 5942, 
    9632, 12412, 18592, 20383, 25453, 26921, 28451, 30589, 31306, 29983, 
    30803, 29210, 27998, 24913, 21136, 19409, 14209, 11236, 6979, 3834, 
    -1560, -4730, -9044, -14177, -17641, -21912, -24050, -26666, -29552, 
    -30188, -30425, -31227, -30598, -29443, -27127, -25767, -22063, -19301, 
    -17069, -10641, -9421, -1988, 1773, 5794, 7765, 15209, 16529, 19446, 
    22889, 25447, 28153, 29025, 30414, 31265, 31089, 28115, 27431, 25470, 
    22968, 19416, 15899, 11465, 9058, 4236, -447, -5039, -10292, -11924, 
    -16689, -21785, -22340, -26588, -28263, -29035, -30017, -30578, -29123, 
    -28162, -27775, -25612, -21481, -18985, -16027, -12387, -7660, -4104, 
    482, 4339, 10758, 13004, 16586, 18767, 22380, 26159, 28715, 28902, 30160, 
    30114, 30593, 29120, 28189, 25242, 21501, 21039, 16102, 13121, 7342, 
    5462, 381, -3497, -9463, -11543, -15438, -20073, -23808, -27288, -27938, 
    -30553, -30241, -32276, -29558, -29933, -29427, -25378, -23688, -20530, 
    -16834, -13106, -8300, -4246, -128, 3243, 7884, 14002, 16903, 21373, 
    24465, 26881, 27132, 29697, 31249, 30689, 29859, 29572, 28297, 26666, 
    24052, 21393, 15587, 13207, 7975, 4830, -1318, -3943, -9027, -12638, 
    -16632, -20299, -23195, -25828, -28835, -30468, -30424, -30890, -30078, 
    -28295, -26423, -26408, -22763, -20456, -18271, -12219, -8540, -4633, 
    -518, 4476, 9594, 11957, 14693, 18913, 21563, 25297, 27828, 30678, 31472, 
    31397, 31125, 29504, 29547, 26157, 23711, 20744, 15348, 13643, 9796, 
    4744, 2024, -4595, -8461, -12176, -15777, -18187, -23800, -25393, -28972, 
    -28615, -31049, -30519, -30163, -29438, -28755, -27935, -23942, -19439, 
    -18612, -15315, -9576, -3630, -538, 4792, 7626, 11976, 15161, 19679, 
    22726, 25819, 26816, 28300, 29564, 30322, 30758, 29523, 28200, 27815, 
    23343, 20894, 17526, 14044, 11316, 5723, 31, -2830, -6482, -10971, 
    -16737, -19573, -23680, -23793, -27566, -28885, -31142, -30880, -29659, 
    -30258, -29781, -26284, -22761, -21260, -17863, -13425, -10823, -5884, 
    -1177, 1406, 6541, 11174, 16657, 19763, 21497, 26545, 26472, 28672, 
    30489, 32091, 30624, 30161, 28567, 25500, 24137, 21118, 18076, 13745, 
    9474, 4772, 301, -2395, -7653, -10925, -14775, -19914, -21777, -25780, 
    -27034, -29911, -30019, -31356, -30285, -29924, -28872, -28151, -23574, 
    -20589, -18535, -15256, -10441, -5729, -2906, 2984, 8133, 9923, 14751, 
    18449, 21642, 25175, 28444, 28437, 30819, 30956, 29530, 30727, 28863, 
    27223, 23360, 21406, 18380, 15272, 11489, 4937, 1632, -1681, -6144, 
    -10838, -15055, -17339, -20627, -24755, -27687, -27905, -31459, -29712, 
    -29851, -30317, -29270, -27445, -23552, -22336, -19125, -13829, -10237, 
    -8001, -2559, 1315, 5062, 8999, 15554, 17549, 21543, 24420, 26075, 28223, 
    30854, 30297, 29761, 31579, 27964, 28480, 25254, 23261, 18892, 13727, 
    11253, 6887, 1753, -1886, -6926, -10445, -14720, -18393, -21789, -25759, 
    -28753, -27757, -30866, -31000, -30563, -31072, -28655, -27333, -24403, 
    -22629, -17815, -15811, -11343, -6577, -2389, 768, 5103, 10169, 15504, 
    18329, 21441, 23340, 27441, 28086, 30661, 30559, 31421, 32011, 29732, 
    27898, 24217, 22249, 20054, 14856, 9921, 7754, 2628, -2099, -4672, -9144, 
    -14592, -19022, -21773, -24280, -25981, -29360, -30149, -31698, -32259, 
    -29031, -27700, -27757, -25121, -21376, -18578, -16881, -10374, -6181, 
    -4010, 2582, 4382, 10414, 13714, 17938, 20477, 25671, 27364, 28326, 
    29566, 30285, 30212, 31540, 29374, 26797, 26392, 23378, 18861, 15670, 
    12734, 7300, 3595, -674, -5910, -9058, -13870, -17120, -22029, -24377, 
    -25304, -28014, -29738, -31530, -30034, -29815, -29384, -29012, -24948, 
    -21696, -18367, -16497, -11620, -7713, -2877, 327, 6766, 9301, 14112, 
    17015, 21032, 24367, 27526, 27860, 29007, 30578, 30270, 30713, 28449, 
    28319, 26050, 22953, 20470, 17656, 11697, 7743, 3768, -983, -5020, -8908, 
    -13102, -15866, -20019, -24290, -27819, -28931, -28883, -32193, -29833, 
    -30753, -29077, -28032, -26824, -22072, -20013, -17563, -12505, -7697, 
    -4604, 143, 3883, 10036, 11548, 17088, 18932, 22553, 26957, 27937, 29103, 
    31290, 31235, 29486, 28025, 28256, 26185, 22981, 20168, 16152, 12522, 
    9225, 3917, -2116, -3476, -9987, -13738, -17808, -20181, -23877, -24969, 
    -27230, -30303, -30693, -29535, -31498, -30380, -26802, -25766, -22589, 
    -20385, -16878, -12884, -7921, -2889, 1624, 3277, 8357, 12397, 17504, 
    20445, 22924, 25627, 29548, 30535, 30604, 32340, 30934, 29118, 26801, 
    25612, 23729, 21819, 16466, 12460, 8654, 5945, 227, -2349, -7114, -12336, 
    -17504, -20143, -22854, -27263, -29255, -29797, -30721, -29713, -31503, 
    -30342, -27676, -26901, -23894, -20389, -15515, -13130, -8070, -6553, 
    -407, 5514, 8162, 13864, 15733, 17915, 22468, 25624, 26450, 30142, 29971, 
    30177, 30895, 30707, 28122, 24982, 23542, 20773, 18393, 14588, 7822, 
    4103, 709, -3093, -9195, -10831, -16016, -18769, -23383, -25441, -27702, 
    -29641, -31130, -31221, -29970, -28503, -27226, -25089, -24680, -19910, 
    -18007, -14669, -8569, -4810, -1008, 2188, 7488, 11955, 14985, 19370, 
    24207, 25992, 26879, 29620, 30792, 29580, 30419, 31133, 27817, 26494, 
    24029, 19399, 15819, 12477, 9330, 6797, 1893, -4910, -7824, -11707, 
    -16469, -18888, -23429, -24055, -25846, -29169, -30490, -31371, -30128, 
    -28644, -28067, -25879, -25505, -21020, -18429, -13230, -10021, -5001, 
    -1786, 2620, 7349, 10909, 15781, 19311, 21238, 24886, 28093, 28172, 
    28654, 30716, 30275, 29045, 29025, 27289, 25036, 20712, 19140, 15148, 
    10119, 5451, 249, -2613, -8525, -11725, -14261, -18831, -22295, -24993, 
    -27264, -29427, -30172, -32233, -30416, -31288, -27855, -26103, -23369, 
    -21948, -18059, -13936, -11189, -4682, -886, 3660, 6445, 10764, 14811, 
    17633, 23047, 25109, 27402, 28314, 28471, 31208, 30763, 31598, 28882, 
    27921, 24964, 21523, 18886, 13269, 10037, 7017, 2743, -2468, -6156, 
    -9755, -14942, -18071, -22706, -25087, -27977, -28605, -30130, -29995, 
    -31705, -30597, -28196, -26083, -26211, -23199, -18246, -15822, -9395, 
    -5033, -2853, 1812, 7087, 9969, 14976, 18589, 21089, 25561, 26843, 27557, 
    31932, 29754, 29138, 29146, 27851, 26702, 24490, 20661, 16918, 14817, 
    10228, 5750, 2137, -1577, -5474, -9236, -13764, -19445, -21759, -23942, 
    -26587, -29611, -29082, -30065, -31377, -31180, -28491, -28695, -25145, 
    -22496, -19623, -16240, -11154, -7270, -3752, 2895, 7001, 11438, 15496, 
    17644, 21894, 23869, 27685, 29056, 30283, 31162, 32064, 31644, 28805, 
    29151, 23967, 22803, 20163, 16128, 11004, 6962, 4269, -806, -5278, -9493, 
    -12579, -18275, -21782, -24468, -27106, -28710, -29037, -31572, -29574, 
    -30397, -28061, -27265, -25475, -23817, -19820, -13822, -10208, -7577, 
    -3960, 2073, 6215, 10572, 13208, 16954, 21408, 24357, 26363, 28441, 
    29667, 29564, 30668, 28754, 29830, 27771, 26178, 22409, 20303, 15203, 
    11209, 7550, 2380, -705, -4389, -9164, -13960, -17230, -20284, -24165, 
    -26744, -27940, -28670, -29835, -32035, -30320, -28724, -27010, -25732, 
    -23595, -19492, -17764, -10797, -8092, -3963, 344, 5672, 10059, 13084, 
    17089, 21578, 24155, 27427, 27385, 31289, 29967, 31468, 31101, 28180, 
    28005, 24989, 22123, 19584, 16782, 10959, 7125, 3428, -1788, -4267, 
    -8204, -13816, -18357, -21797, -22480, -25538, -28613, -30774, -30999, 
    -30102, -30719, -30126, -28059, -26328, -24608, -19055, -16762, -12506, 
    -8926, -4528, 1073, 3418, 10814, 14949, 17936, 21190, 22136, 24930, 
    27226, 30509, 30493, 32411, 31351, 29587, 27052, 26562, 23515, 19245, 
    17455, 11961, 8934, 3381, 512, -4303, -8409, -13962, -15591, -19085, 
    -22775, -26776, -27229, -28816, -30202, -31734, -30340, -29404, -28425, 
    -25131, -23145, -19846, -18433, -13102, -8465, -5397, 248, 5857, 8314, 
    13304, 17205, 21795, 21554, 26040, 27970, 31014, 29373, 31430, 30903, 
    27927, 27185, 25382, 23129, 19103, 17541, 13459, 8639, 4789, 990, -3457, 
    -8611, -11832, -16912, -19554, -21208, -26225, -29362, -28982, -29115, 
    -30830, -30575, -31072, -27443, -27092, -23877, -21850, -15327, -11876, 
    -9963, -4505, -460, 3534, 7838, 12238, 16223, 19505, 22456, 25638, 28712, 
    29342, 29512, 30670, 31084, 29114, 29143, 26437, 23628, 20542, 16904, 
    13527, 9826, 4710, 418, -2350, -8111, -12064, -16448, -19665, -23299, 
    -25166, -27120, -29921, -30652, -29496, -31878, -30193, -29714, -27161, 
    -24114, -19984, -17545, -13432, -9203, -5409, -542, 4725, 8159, 10667, 
    15491, 19661, 23344, 25082, 27610, 28086, 28975, 30478, 29708, 29781, 
    26984, 26109, 24993, 21248, 18067, 13757, 9859, 5480, -595, -3938, -6736, 
    -11375, -15664, -18701, -22104, -26447, -27609, -28273, -30253, -31653, 
    -30649, -31006, -28136, -26740, -23796, -22240, -17788, -14516, -9849, 
    -5817, -2149, 2496, 8046, 12382, 15636, 17940, 22336, 25238, 29105, 
    29155, 30416, 30696, 30749, 30490, 29671, 25597, 23025, 21112, 17176, 
    13753, 10536, 5544, 1522, -2981, -5368, -11100, -15870, -19427, -23536, 
    -25161, -27474, -30483, -31010, -31297, -32149, -29104, -28245, -27288, 
    -24349, -21675, -19109, -12660, -10124, -6002, -421, 1472, 6471, 12278, 
    13950, 19895, 21752, 24861, 27377, 28513, 30579, 31469, 32142, 28999, 
    27725, 26391, 24845, 21826, 19746, 14844, 10745, 5380, 2333, -1266, 
    -6959, -10807, -15107, -19515, -21620, -25100, -26787, -30139, -30097, 
    -30421, -30878, -31052, -28341, -28294, -24085, -21349, -18426, -15362, 
    -11364, -8000, -3457, 1422, 6200, 11236, 14065, 17194, 22466, 24319, 
    26204, 29856, 30706, 31623, 30610, 30536, 29395, 27186, 25045, 22089, 
    18996, 15551, 12254, 7076, 3183, -3894, -6373, -10167, -13303, -17037, 
    -22840, -24582, -25941, -28547, -30966, -30161, -30289, -29765, -29253, 
    -27700, -23862, -22837, -19703, -14729, -11507, -5576, -2241, 1692, 5251, 
    11117, 13765, 17837, 21674, 24923, 27272, 28662, 28961, 30433, 29860, 
    30395, 30231, 26141, 24096, 22070, 20338, 16274, 11400, 7611, 3142, 
    -2439, -5983, -11310, -14009, -16485, -20432, -24156, -26904, -28579, 
    -28808, -30262, -31906, -30915, -29034, -28614, -25412, -22999, -18426, 
    -15100, -10712, -7710, -3227, 1276, 5344, 9231, 13678, 17559, 21848, 
    23920, 25737, 28770, 29853, 30859, 30837, 31007, 28844, 28490, 26853, 
    23474, 18742, 15723, 11688, 7187, 2118, -1355, -4538, -8046, -13031, 
    -17747, -21636, -23114, -25252, -27061, -29566, -28982, -30752, -29288, 
    -29812, -27097, -26288, -22885, -17703, -14508, -13611, -6215, -3131, 
    371, 4334, 9842, 11893, 17404, 19756, 24525, 26714, 29360, 29861, 30638, 
    31179, 29395, 30493, 26451, 26963, 23303, 18361, 16588, 12556, 9304, 
    3481, -167, -5956, -10588, -12811, -17255, -21018, -24290, -26000, 
    -27103, -30527, -29354, -30704, -30334, -29581, -27634, -26962, -23531, 
    -19550, -15784, -12571, -7964, -3069, -543, 5629, 9915, 11684, 15530, 
    20251, 24079, 26279, 28893, 29777, 30376, 31987, 31321, 28824, 27238, 
    25759, 22681, 18645, 17105, 11287, 8697, 4542, -1399, -3336, -8529, 
    -12026, -15436, -20930, -23760, -26898, -27553, -28637, -30336, -31171, 
    -29438, -30015, -27990, -24787, -22241, -20574, -14808, -14238, -9312, 
    -5667, 1817, 3822, 7676, 13204, 16041, 20451, 23133, 26966, 28602, 29075, 
    31434, 32418, 30008, 27926, 28126, 25423, 23526, 19395, 17693, 14123, 
    9863, 4041, 411, -4268, -8200, -13155, -16879, -19396, -22445, -25500, 
    -26585, -29294, -30164, -31757, -30547, -29218, -27883, -27902, -22958, 
    -19781, -16478, -14066, -7922, -4933, 6, 2861, 6840, 12478, 15940, 18670, 
    22356, 25580, 27709, 29504, 31388, 31601, 29031, 28941, 27927, 27477, 
    22795, 21446, 17389, 11939, 10142, 5265, 111, -4152, -8281, -11121, 
    -17381, -19888, -22629, -24819, -27696, -28405, -30147, -29639, -30313, 
    -30530, -28425, -24892, -23799, -21062, -16163, -14090, -11193, -5714, 
    698, 4575, 8655, 13487, 14922, 18997, 22849, 25788, 27868, 30437, 30670, 
    31978, 31714, 29746, 28293, 26906, 25680, 21031, 17565, 13717, 9502, 
    7007, -284, -2773, -8971, -11550, -14812, -20185, -23018, -25826, -26732, 
    -27993, -29250, -31025, -29912, -30422, -28155, -26884, -22557, -20595, 
    -16641, -14002, -10189, -6745, -1458, 2578, 7367, 12586, 16907, 19826, 
    22106, 26884, 27413, 27602, 30939, 30524, 31978, 30040, 28692, 27176, 
    23336, 21160, 17393, 15407, 10138, 5697, 2423, -3852, -8015, -12593, 
    -14619, -19229, -22071, -24350, -28603, -28945, -30821, -32006, -31815, 
    -30191, -29286, -26524, -24657, -21967, -18298, -14330, -10413, -5555, 
    -1917, 2851, 6579, 11581, 13600, 19405, 23063, 25701, 28722, 28825, 
    31023, 30836, 29946, 30064, 28660, 25616, 24534, 21122, 18525, 14938, 
    11676, 6799, 2249, -3433, -6951, -10561, -14443, -18625, -21815, -23983, 
    -25572, -28148, -28425, -30999, -31203, -28733, -28870, -27409, -24362, 
    -22599, -19537, -14317, -10602, -5794, -3638, 3059, 7893, 10867, 14200, 
    18936, 21308, 23851, 27603, 30430, 30162, 31441, 31565, 30804, 29585, 
    25513, 24645, 23004, 19596, 15093, 11755, 6525, 4251, -2077, -8115, 
    -9937, -14504, -16856, -20468, -24238, -26574, -27762, -29091, -30001, 
    -31202, -29382, -27969, -27391, -25352, -22062, -19635, -14149, -11148, 
    -7569, -3903, 2464, 6869, 11822, 14387, 17445, 20940, 24761, 27462, 
    30060, 28809, 31084, 30182, 29820, 28221, 28298, 24659, 22163, 19933, 
    14234, 11911, 8074, 1544, -1989, -6308, -10540, -14828, -17591, -21119, 
    -24720, -26774, -29440, -30395, -30509, -31394, -29754, -29626, -25651, 
    -26803, -23093, -18149, -15717, -11355, -6027, -2972, 1633, 5978, 8989, 
    13392, 17792, 20807, 22446, 27719, 29311, 30888, 31604, 30456, 30183, 
    29153, 27179, 24466, 22497, 20852, 15965, 11349, 8222, 2329, -749, -6211, 
    -8785, -13006, -17090, -21452, -23947, -26202, -29020, -29137, -31856, 
    -30395, -29559, -27617, -28339, -25490, -23378, -18760, -16119, -13001, 
    -7924, -3536, 1666, 5679, 8971, 13116, 18626, 21624, 24802, 25335, 28092, 
    30028, 30592, 30930, 31440, 29573, 27507, 25359, 22054, 18684, 15005, 
    13824, 6758, 3979, -1076, -3355, -9149, -14075, -17381, -21429, -22569, 
    -25533, -27274, -28549, -30058, -30903, -31154, -28726, -29430, -24220, 
    -21423, -19946, -17177, -12734, -7854, -4800, 993, 4745, 9987, 12852, 
    17486, 20935, 21965, 25589, 28226, 30288, 31071, 31396, 31761, 30767, 
    27773, 24274, 23440, 20647, 17545, 12646, 7645, 3559, -1646, -4465, 
    -8909, -13671, -18518, -19833, -23153, -26282, -27505, -28497, -28771, 
    -31586, -30821, -28864, -28982, -27140, -22935, -19763, -17935, -12446, 
    -7738, -2896, -537, 3980, 8135, 13240, 17313, 21231, 24168, 25128, 28790, 
    29466, 29307, 30064, 31533, 29693, 27355, 26996, 22358, 21350, 16421, 
    12139, 9983, 3981, 1899, -3557, -8638, -12777, -17179, -20975, -22718, 
    -25592, -27841, -29793, -31343, -31156, -31934, -28529, -26626, -25812, 
    -24323, -21136, -17410, -14579, -7640, -5391, -21, 5572, 9017, 11998, 
    16942, 20040, 23309, 25675, 26797, 31081, 29323, 29935, 28702, 29502, 
    27904, 25873, 22860, 21588, 16340, 13623, 10168, 6056, -95, -3254, -9573, 
    -11571, -15450, -20542, -23211, -25173, -27579, -29243, -31363, -30942, 
    -31414, -29340, -29145, -26584, -23937, -20093, -17755, -12080, -8719, 
    -5442, -27, 4166, 7763, 10763, 14688, 19004, 22068, 25819, 27117, 30611, 
    31698, 31123, 29168, 30134, 28461, 27592, 22968, 19411, 17795, 12585, 
    9348, 5904, 1681, -3537, -7593, -11550, -16506, -19118, -21110, -25136, 
    -26263, -28814, -28995, -32163, -29967, -31049, -29382, -25988, -24046, 
    -19796, -18265, -13850, -8908, -5059, -2085, 4696, 7457, 9851, 15355, 
    18854, 21696, 24026, 26625, 30370, 29623, 30436, 29499, 30110, 29775, 
    26045, 25085, 20175, 16050, 14774, 8799, 7417, 1938, -2631, -7105, 
    -12272, -14932, -20650, -22782, -26119, -27138, -27774, -30297, -31705, 
    -31152, -30968, -28394, -27425, -23605, -21724, -17592, -14289, -10729, 
    -5794, -668, 2762, 5965, 12213, 15361, 19727, 22961, 25017, 27048, 28664, 
    29748, 30199, 30233, 29743, 28426, 27186, 24522, 20820, 19071, 14910, 
    10572, 7024, 1158, -2277, -8220, -10571, -14747, -19749, -21438, -24093, 
    -25527, -28947, -29526, -30078, -31244, -31674, -28932, -27226, -25093, 
    -21204, -18410, -15811, -12112, -5740, -965, 1479, 7556, 9406, 14607, 
    19050, 20744, 24306, 27864, 29825, 29794, 31041, 31243, 30016, 29907, 
    26756, 24760, 22824, 20275, 15698, 9941, 7137, 4075, -1834, -6065, -9949, 
    -14877, -18603, -21234, -25121, -26857, -27934, -30803, -30112, -28971, 
    -31699, -27482, -26505, -24360, -22905, -17016, -14934, -11296, -6756, 
    -2174, 2569, 6820, 9871, 14243, 18676, 21491, 23330, 26506, 28496, 30645, 
    30029, 32386, 30959, 28158, 26393, 25014, 21348, 19367, 15292, 10646, 
    7724, 2152, -2559, -6142, -9084, -14539, -19145, -21046, -25589, -28237, 
    -30052, -29459, -30332, -31898, -30317, -30089, -27902, -24286, -21805, 
    -20621, -16039, -10277, -6609, -2628, 832, 7090, 10331, 13940, 17892, 
    21299, 24670, 27785, 28413, 28535, 29973, 29842, 29526, 29338, 27876, 
    24805, 23041, 19395, 15602, 12473, 9052, 4139, -747, -5168, -10245, 
    -13291, -17618, -22040, -24045, -25802, -28872, -30787, -30456, -32164, 
    -30858, -29816, -27017, -25573, -21568, -18486, -16479, -10967, -9104, 
    -3507, 1491, 5327, 9468, 12586, 15705, 20458, 22902, 27569, 27660, 30058, 
    30761, 31356, 30613, 28458, 28826, 26101, 22559, 19399, 14618, 11926, 
    8119, 3962, -761, -5465, -8793, -13512, -17145, -22128, -23795, -26403, 
    -28017, -28461, -29641, -31315, -30935, -29381, -27642, -25837, -22337, 
    -19629, -15498, -13778, -7490, -3287, 96, 5684, 9469, 12368, 16488, 
    19987, 22148, 27076, 28705, 29786, 29911, 30208, 30364, 30222, 29593, 
    25249, 23283, 20213, 15710, 14095, 8211, 4476, -1358, -4556, -8385, 
    -11689, -17437, -18691, -22372, -26783, -28439, -30087, -30996, -32573, 
    -30605, -29305, -28313, -24998, -22592, -19093, -15840, -12810, -9159, 
    -4339, 806, 5368, 7341, 12641, 15729, 19655, 24025, 25290, 26577, 28178, 
    30435, 31159, 30104, 28579, 27976, 25817, 22581, 20032, 17011, 12915, 
    8523, 5776, 12, -4683, -9501, -13532, -16667, -19556, -22882, -26231, 
    -27874, -28841, -31083, -29709, -31334, -30125, -28794, -25315, -23453, 
    -19138, -16161, -14860, -8364, -4487, -757, 3347, 9089, 11117, 16393, 
    19397, 22840, 26452, 27642, 29613, 30700, 31210, 32272, 30484, 27081, 
    25659, 23782, 19233, 15875, 11792, 8858, 4653, 498, -5327, -8139, -12645, 
    -15764, -19475, -22523, -26155, -28531, -29971, -31241, -31376, -31552, 
    -29302, -29283, -26088, -23738, -21741, -17495, -14172, -9953, -4562, 
    -206, 2718, 8410, 12304, 15614, 20229, 23665, 25678, 27095, 30191, 31311, 
    30976, 32008, 28643, 27134, 24898, 22411, 20815, 16716, 12613, 9941, 
    5240, 2098, -2026, -8623, -12430, -17375, -19850, -22932, -24298, -27777, 
    -29243, -29993, -31525, -30449, -30255, -28143, -26635, -23296, -21609, 
    -18578, -12433, -10827, -4826, -2520, 2906, 7657, 12167, 14269, 18869, 
    21021, 25191, 28697, 30309, 31785, 31975, 31555, 30137, 28474, 27569, 
    24971, 20631, 18952, 13998, 9368, 5850, 95, -3201, -7728, -9612, -15572, 
    -19781, -23570, -24982, -26825, -28769, -29523, -30819, -30345, -30480, 
    -27897, -27775, -24867, -22987, -17464, -13946, -11041, -5738, -1811, 
    3004, 7237, 11440, 16310, 19344, 21794, 24803, 27134, 27343, 30626, 
    31467, 30852, 30132, 28223, 25311, 24475, 20467, 18030, 14907, 10669, 
    6696, 2076, -2742, -6519, -11296, -15219, -19292, -21390, -26521, -26273, 
    -29996, -29038, -31343, -31745, -31581, -30054, -27995, -24781, -21957, 
    -19458, -15467, -11781, -7261, -2377, 770, 8098, 10962, 15970, 16912, 
    22961, 25511, 26790, 29198, 30750, 30442, 29333, 29821, 30087, 27188, 
    24095, 23137, 19615, 13857, 12453, 5493, 3709, -1664, -7108, -11680, 
    -14890, -17161, -22673, -24669, -26028, -27214, -30287, -31785, -30838, 
    -30316, -30417, -27874, -25511, -22283, -20301, -15985, -11894, -6738, 
    -3336, 829, 5993, 8476, 15575, 18433, 19920, 24834, 27007, 28515, 28864, 
    31372, 31080, 30541, 28387, 26863, 25327, 23201, 20220, 15445, 12610, 
    6132, 2923, -1127, -6024, -10098, -13590, -17067, -20354, -24332, -25718, 
    -28724, -29948, -30891, -31078, -31518, -30423, -27198, -25396, -20647, 
    -18941, -15294, -12657, -8888, -3142, 1028, 4667, 8547, 13711, 17527, 
    22129, 23332, 26287, 28859, 29639, 31618, 32040, 29356, 28555, 27555, 
    23455, 22474, 18457, 16930, 12038, 7476, 3854, 205, -5550, -8124, -12144, 
    -18620, -22374, -22596, -27538, -27970, -30000, -31379, -29993, -30405, 
    -29537, -26481, -24392, -21493, -19186, -16957, -11409, -7147, -4634, 
    1625, 5239, 8665, 12345, 17868, 19638, 22859, 26016, 29614, 30231, 29938, 
    30052, 31643, 28252, 27680, 25852, 23657, 18028, 15730, 12037, 7202, 
    4793, 526, -4176, -9156, -13121, -16704, -20260, -25303, -27899, -29592, 
    -31087, -30776, -29801, -30365, -29795, -27001, -24487, -23240, -18182, 
    -16216, -13105, -8247, -4988, 380, 4828, 8188, 13754, 17086, 21074, 
    22379, 25925, 27881, 29602, 30572, 30518, 30156, 29107, 27350, 25077, 
    23493, 18578, 16412, 13185, 9034, 3096, -1510, -5028, -8721, -13463, 
    -16806, -20394, -23280, -27087, -29297, -30265, -30193, -31007, -32071, 
    -31112, -29391, -24763, -24395, -20695, -17511, -13261, -8704, -3656, 
    773, 4397, 9027, 13047, 15483, 21166, 24979, 26829, 27662, 29548, 31295, 
    32139, 30245, 28530, 28585, 25929, 22928, 19644, 15830, 13696, 8125, 
    5486, 194, -3398, -8636, -11209, -17826, -19397, -21548, -25773, -27269, 
    -28922, -30007, -32343, -30839, -30951, -28814, -26666, -22387, -20798, 
    -17540, -14386, -8704, -4975, 288, 4467, 8066, 11635, 16470, 18299, 
    22991, 27072, 29126, 29445, 30412, 31612, 31840, 30489, 29177, 25356, 
    23173, 20253, 16932, 13149, 8997, 4799, 461, -3917, -8284, -12727, 
    -16734, -20814, -24294, -23970, -28461, -29567, -31844, -29221, -30053, 
    -30339, -28149, -26153, -22601, -20999, -15970, -13755, -8996, -5681, 
    -383, 2254, 8540, 12656, 14852, 19948, 23469, 24297, 27109, 30213, 31334, 
    29773, 30356, 30506, 29697, 26862, 23229, 21915, 16806, 11837, 9936, 
    4837, 494, -3232, -8080, -13180, -15658, -19249, -22292, -26301, -27817, 
    -29180, -31335, -30183, -29789, -30624, -28301, -27712, -24569, -22676, 
    -16964, -15009, -10206, -4325, -2264, 3923, 7599, 12085, 15740, 18455, 
    22617, 26448, 26615, 28065, 29169, 31433, 30768, 29350, 28359, 27214, 
    24710, 21405, 19508, 13514, 10239, 5867, 1771, -2324, -7557, -10552, 
    -15863, -19970, -23554, -24437, -27080, -28616, -30806, -29123, -29522, 
    -28778, -26799, -27760, -24219, -20918, -17554, -13001, -10695, -7269, 
    -1809, 1316, 6704, 10716, 14099, 18802, 22530, 25381, 26731, 29161, 
    29861, 29182, 30046, 30684, 28970, 27960, 24492, 22505, 17313, 14046, 
    11139, 5187, 1390, -3749, -7853, -10431, -16092, -20124, -22283, -24704, 
    -26827, -28889, -31050, -30493, -31342, -30692, -28524, -27694, -26285, 
    -21195, -17880, -14131, -10735, -7948, -2612, 2649, 7935, 10086, 14614, 
    17298, 20190, 24377, 25443, 28800, 29994, 31400, 30249, 30438, 28999, 
    26971, 24403, 21988, 20069, 14857, 10421, 6920, 2453, -1616, -6894, 
    -11836, -15281, -17644, -20776, -23727, -26752, -27920, -29437, -32202, 
    -31977, -29964, -29725, -26031, -26157, -23500, -18347, -14417, -11343, 
    -7458, -2346, 2472, 5940, 9900, 14167, 18681, 21287, 24377, 25919, 27040, 
    29127, 31473, 31665, 30996, 30452, 27048, 24845, 22320, 19916, 14501, 
    10142, 7995, 2623, -1168, -6723, -11037, -13825, -18722, -22677, -23405, 
    -26433, -27534, -30157, -30413, -30855, -29919, -27779, -28541, -25218, 
    -22516, -19156, -14952, -11648, -6452, -3480, 1641, 6589, 10770, 14897, 
    17706, 20486, 23330, 24780, 28283, 29994, 30956, 31306, 31536, 28901, 
    28445, 25735, 22522, 19677, 17235, 12214, 6968, 3538, -29, -5780, -9733, 
    -13373, -18513, -20872, -25011, -26615, -27288, -29697, -30632, -30877, 
    -29211, -29501, -27768, -25304, -21870, -18427, -14546, -10646, -7263, 
    -3130, 1594, 6275, 8709, 15417, 17224, 22041, 24769, 27136, 26782, 30441, 
    31142, 30653, 29575, 29226, 26770, 24992, 22111, 19917, 15850, 11565, 
    8479, 2266, -976, -5253, -8175, -15186, -17370, -20849, -23772, -27040, 
    -26593, -30001, -30151, -29970, -31223, -30778, -27726, -25595, -23610, 
    -20490, -16457, -11367, -8710, -2829, 34, 5723, 10501, 13195, 18517, 
    19086, 22584, 26122, 28572, 30424, 29983, 31219, 29787, 29781, 27879, 
    24321, 22645, 21109, 16773, 12119, 7775, 3650, 20, -4279, -8489, -13121, 
    -16118, -19865, -23362, -24818, -27303, -28792, -30108, -30593, -30621, 
    -29737, -28281, -25813, -22065, -21365, -16157, -11933, -9196, -3207, 
    -250, 5809, 7793, 12278, 15068, 21051, 22231, 26665, 28236, 28812, 30183, 
    29652, 30954, 29389, 27299, 26750, 22943, 21383, 16084, 13139, 7779, 
    4960, 38, -5323, -8777, -12395, -15761, -21558, -23686, -26847, -27087, 
    -29839, -30564, -30314, -31499, -28730, -29442, -27975, -23430, -19979, 
    -16822, -12660, -8322, -5036, -527, 4849, 8996, 11115, 16942, 20331, 
    22590, 26006, 27916, 29403, 31248, 29841, 31887, 29974, 28042, 25879, 
    23528, 21586, 15875, 12601, 8510, 5323, 2155, -4508, -7406, -13835, 
    -15691, -19957, -22752, -25808, -26883, -28403, -29929, -30366, -31039, 
    -29037, -28376, -26954, -23117, -22091, -18056, -13897, -10948, -4879, 
    -226, 3157, 8496, 13175, 16337, 18720, 22601, 26767, 28660, 28992, 30794, 
    31198, 30999, 30928, 28771, 25770, 22816, 20144, 16798, 13938, 9545, 
    4940, 694, -3806, -7796, -10282, -16296, -18972, -22895, -25242, -29110, 
    -28303, -30723, -29119, -30834, -29944, -28563, -26816, -22422, -21402, 
    -18753, -14390, -10349, -4862, -1230, 3258, 5936, 11863, 16843, 20322, 
    23521, 26219, 27083, 28238, 29217, 32027, 29314, 28814, 28989, 25339, 
    24485, 21017, 17887, 12880, 10135, 5771, 2926, -2349, -6192, -12626, 
    -14255, -19310, -21974, -26227, -26681, -30298, -30272, -31609, -31240, 
    -30236, -29997, -26518, -24339, -21945, -18470, -13990, -10735, -5440, 
    -2939, 1812, 7503, 11849, 13573, 18150, 20992, 24500, 27108, 28471, 
    30033, 30439, 31008, 30210, 27886, 27558, 24914, 21770, 19798, 12950, 
    10708, 5917, 1700, -1807, -7141, -12198, -13888, -17561, -22516, -24267, 
    -27443, -28733, -29372, -30390, -30078, -30198, -29602, -27493, -25931, 
    -22088, -19289, -14911, -9441, -6398, -1716, 2447, 5342, 11025, 15604, 
    19081, 21869, 24564, 27893, 28005, 29978, 30630, 29904, 29055, 28556, 
    26761, 25405, 22500, 19791, 15228, 11992, 7088, 1990, -2547, -6411, 
    -9726, -15663, -19347, -21923, -24153, -26666, -30039, -29786, -31575, 
    -29608, -30193, -29899, -26163, -24835, -22364, -20408, -15713, -10696, 
    -6420, -4408, 2853, 5107, 9238, 13496, 17847, 19767, 23875, 26831, 29616, 
    30025, 31175, 30417, 30182, 28107, 26591, 26432, 20686, 19805, 15376, 
    11681, 8004, 2272, -2228, -5484, -9802, -12959, -18008, -20665, -24232, 
    -26628, -28984, -30276, -30829, -30371, -29744, -30670, -26368, -24274, 
    -22121, -20969, -15464, -10730, -8969, -3490, 2728, 6332, 10640, 14338, 
    19072, 20641, 25057, 25934, 28110, 30352, 30317, 31133, 31531, 28667, 
    28283, 25281, 21127, 18536, 15750, 12291, 8963, 4558, -701, -5174, -9975, 
    -14579, -18432, -21223, -24447, -25625, -28140, -28968, -30656, -31366, 
    -29024, -28881, -27030, -26911, -22465, -19505, -14529, -12522, -9206, 
    -3234, -378, 5693, 8123, 14155, 18046, 19304, 24667, 26078, 28500, 30667, 
    30786, 29233, 31146, 30425, 26243, 24884, 22020, 18544, 15631, 11021, 
    8159, 2565, -1512, -3595, -7863, -13350, -16719, -19754, -23249, -26868, 
    -28709, -30067, -30993, -30694, -28921, -28817, -27786, -25299, -21942, 
    -19690, -15816, -11861, -8610, -5542, 1756, 3618, 8034, 12538, 15984, 
    20142, 22871, 26598, 28709, 28093, 30536, 30313, 31755, 29993, 28419, 
    24650, 23926, 19293, 16523, 12481, 7217, 4388, -290, -4363, -8709, 
    -13481, -17213, -21570, -22718, -26514, -27644, -29696, -29952, -30595, 
    -31558, -29366, -27331, -25859, -22421, -21031, -16812, -13083, -8717, 
    -4022, -435, 4620, 7787, 13212, 17299, 20434, 24858, 26329, 27055, 28178, 
    32392, 30462, 31237, 29967, 27591, 26381, 24609, 21349, 17257, 11742, 
    8475, 4146, -820, -5811, -8200, -13733, -17006, -20163, -22558, -25490, 
    -28876, -29428, -30939, -29342, -29642, -29284, -28072, -24749, -23783, 
    -19769, -17651, -12213, -7270, -5805, 861, 3531, 7963, 12456, 16702, 
    18445, 22316, 26123, 27307, 30147, 31869, 30921, 30122, 28555, 28516, 
    26078, 23126, 20391, 16366, 11913, 7900, 3695, -517, -2382, -8768, 
    -12446, -16192, -19479, -24260, -26260, -27807, -30852, -30780, -29195, 
    -31307, -29071, -27679, -25034, -23001, -19968, -17983, -13662, -10420, 
    -5209, -537, 4259, 6437, 12289, 16860, 19088, 23052, 26966, 27714, 29176, 
    31713, 30874, 30800, 30087, 27977, 26664, 23426, 20154, 17872, 14019, 
    10823, 6611, 298, -3986, -7268, -11109, -14987, -17816, -24107, -26180, 
    -27391, -28711, -29727, -29268, -30993, -31380, -28611, -27146, -23417, 
    -19849, -16314, -14360, -10411, -4564, -2259, 3135, 7558, 9861, 16474, 
    19663, 23710, 23750, 27024, 27877, 30660, 29464, 30449, 29804, 27376, 
    26869, 23854, 21580, 17158, 14151, 10285, 5884, 294, -3373, -6417, 
    -10629, -15244, -19398, -22205, -24974, -27493, -27824, -30300, -30560, 
    -31357, -30248, -28669, -25637, -25067, -21907, -17566, -13636, -10408, 
    -6366, -2424, 2804, 5589, 9688, 15323, 18448, 22864, 23805, 28083, 29808, 
    29238, 29268, 30932, 31175, 27318, 27148, 25613, 21188, 17427, 15691, 
    9566, 6106, 2434, -4235, -7332, -10055, -14656, -19245, -22291, -24881, 
    -26388, -29406, -30764, -31754, -30696, -29972, -29561, -27821, -25219, 
    -20198, -17820, -13872, -10950, -7847, -3317, 2368, 6522, 12037, 14944, 
    18885, 21932, 26089, 27348, 30580, 29229, 31523, 30748, 29686, 29541, 
    27322, 25187, 22571, 18498, 13848, 11231, 6292, 3229, -3148, -6398, 
    -9645, -13128, -17672, -22295, -23541, -28586, -29529, -30761, -29373, 
    -30273, -29481, -30382, -26236, -25209, -21172, -18705, -13874, -10463, 
    -7710, -1979, 2546, 6657, 8661, 13011, 17771, 21735, 25143, 27237, 29819, 
    28761, 30844, 32023, 29214, 28584, 27629, 25707, 22138, 18684, 14674, 
    11477, 5548, 2912, -1164, -6259, -10566, -13787, -17779, -20956, -22918, 
    -25920, -27809, -31606, -30109, -30473, -30525, -29358, -26027, -26130, 
    -22205, -18926, -14374, -10171, -7506, -2621, 652, 5670, 9089, 14694, 
    18199, 20503, 24289, 26589, 29060, 28585, 30863, 29537, 30664, 30223, 
    27339, 26468, 21581, 18177, 14738, 11515, 6299, 3442, -335, -5897, -9207, 
    -12828, -17607, -21015, -25074, -25779, -28766, -29281, -30562, -31339, 
    -30796, -29964, -28108, -24974, -21732, -19910, -16259, -11726, -7676, 
    -4296, 634, 5609, 10111, 12458, 18707, 21131, 23077, 26228, 29158, 30083, 
    30199, 32299, 29873, 28579, 26773, 25551, 24302, 17994, 15289, 12907, 
    9271, 4076, -714, -4810, -9518, -13167, -16378, -21253, -22636, -25399, 
    -28157, -31246, -30552, -31646, -31134, -30049, -28347, -26836, -22081, 
    -20255, -15397, -11399, -7949, -4583, 1247, 5484, 9437, 13954, 15534, 
    20424, 23669, 26231, 29139, 28910, 31288, 30216, 30549, 29394, 28844, 
    25847, 23591, 20452, 16503, 12419, 7974, 4252, 194, -3781, -8577, -13302, 
    -17331, -20659, -24701, -25521, -28934, -30972, -29375, -30402, -29636, 
    -28913, -26983, -26492, -23091, -20394, -17366, -12289, -8254, -3757, 
    1230, 5122, 9193, 13061, 16061, 19271, 23153, 24668, 28470, 29511, 31237, 
    32197, 29542, 30075, 28434, 27008, 23347, 19379, 17075, 13876, 7968, 
    5969, -249, -4209, -7955, -12228, -15496, -21152, -23002, -27020, -28526, 
    -29621, -30356, -30782, -29815, -30999, -28770, -25450, -22024, -21917, 
    -15782, -11734, -8149, -5578, 103, 4636, 7243, 12924, 16790, 20648, 
    22836, 25588, 26885, 28092, 31589, 29897, 30756, 28384, 28507, 26599, 
    25281, 20979, 17206, 14273, 8730, 5964, -516, -3998, -8031, -12873, 
    -15121, -19124, -22688, -26106, -26064, -30967, -30327, -30942, -29861, 
    -30641, -28100, -26161, -25648, -21536, -17698, -12524, -8686, -4925, 
    -1508, 3397, 7463, 11567, 15784, 19371, 23472, 25108, 27628, 30051, 
    30174, 29018, 31381, 30652, 28525, 26628, 25348, 19481, 17228, 12720, 
    10271, 6846, 298, -3708, -8661, -12440, -16467, -18844, -23036, -25536, 
    -28124, -29077, -30959, -30866, -29836, -28382, -29574, -26737, -23908, 
    -21093, -17080, -15186, -10885, -5113, -2031, 2435, 8170, 10363, 14959, 
    18571, 21929, 26195, 28533, 28066, 29906, 29591, 29020, 30364, 27931, 
    25950, 23296, 20902, 17673, 13063, 9588, 6356, 1097, -3420, -8364, 
    -10695, -16710, -19143, -22016, -24950, -27767, -27530, -31169, -31925, 
    -29663, -30287, -30183, -27773, -24367, -20562, -17304, -14609, -8852, 
    -6509, -1558, 2430, 7533, 12277, 14063, 18476, 22937, 25747, 28173, 
    30241, 29635, 31017, 32196, 30945, 27181, 27777, 25899, 21636, 18862, 
    14365, 10197, 7529, 2758, -2061, -7895, -11002, -15204, -20025, -23244, 
    -23335, -26806, -29999, -29705, -29147, -31475, -30258, -29199, -26095, 
    -24904, -21250, -19180, -16627, -10595, -7298, -2971, 3193, 6559, 11862, 
    13925, 18298, 21178, 24503, 27643, 29440, 30051, 30825, 29596, 29183, 
    28324, 27220, 26390, 23453, 18077, 14509, 11776, 5048, 1873, -1092, 
    -6524, -10147, -15354, -18085, -22062, -23941, -27477, -29352, -30181, 
    -31191, -30795, -29761, -28828, -28406, -23851, -21718, -19186, -16193, 
    -10739, -6706, -1920, 2651, 5780, 10038, 15308, 17663, 19820, 24811, 
    26017, 30460, 31342, 30683, 30696, 29298, 29234, 27534, 24205, 22773, 
    17881, 15251, 10959, 8020, 1525, -908, -6573, -10067, -13364, -17984, 
    -21256, -24116, -26526, -28367, -31026, -32206, -31521, -30816, -29519, 
    -28490, -24774, -23889, -17879, -14916, -12318, -6731, -2521, 1163, 5321, 
    8940, 13405, 17513, 21372, 24028, 26976, 28112, 30339, 30292, 30142, 
    31217, 29033, 26708, 24817, 22773, 18437, 17072, 11380, 7877, 4077, 326, 
    -4842, -10583, -12730, -17179, -21990, -23124, -25346, -27850, -29559, 
    -30818, -30306, -29496, -29636, -27672, -24247, -22180, -19104, -15761, 
    -12121, -8556, -2473, -459, 6438, 8228, 13205, 16691, 19992, 24918, 
    25535, 27591, 28855, 30486, 29926, 31988, 29147, 26886, 25492, 21665, 
    19021, 17433, 11838, 7967, 5409, -2351, -5889, -10435, -13974, -18372, 
    -19115, -24633, -26972, -28890, -28456, -30199, -30567, -29323, -29526, 
    -26596, -25382, -22234, -19946, -16299, -13727, -7478, -3916, 455, 4789, 
    8690, 13318, 17693, 20486, 24184, 25362, 29360, 29886, 31988, 29981, 
    30599, 29972, 27776, 25795, 23841, 19093, 16318, 13434, 7954, 4231, 
    -1075, -4715, -8776, -12615, -15207, -20283, -24104, -25819, -29726, 
    -29117, -30795, -31725, -31848, -30224, -27226, -26584, -23241, -20623, 
    -16027, -13840, -9727, -5325, 1594, 4596, 9516, 12580, 16442, 19946, 
    23851, 24512, 27164, 31358, 29762, 31919, 30361, 29004, 27323, 25974, 
    23300, 18841, 17398, 12577, 9117, 3132, 1239, -2953, -9113, -13185, 
    -15403, -20846, -21979, -25077, -27019, -29414, -29422, -30581, -31583, 
    -30693, -27525, -26324, -24056, -19306, -18376, -12406, -8950, -3635, 
    -1956, 3186, 8992, 12337, 14869, 18019, 22705, 25966, 28880, 29116, 
    30222, 32528, 29139, 30165, 27746, 26789, 23520, 21207, 17063, 12981, 
    9460, 3310, -144, -4179, -8161, -12631, -17722, -20068, -23715, -25480, 
    -27321, -29674, -30476, -30965, -30884, -29463, -28329, -26471, -23974, 
    -21033, -17615, -13506, -9809, -4602, -2219, 2228, 8574, 12384, 15513, 
    18926, 22818, 24330, 28290, 29164, 31026, 30415, 30487, 29273, 29397, 
    26922, 25763, 21759, 18213, 13835, 9960, 4648, 528, -3888, -8548, -11427, 
    -16624, -18362, -22824, -26187, -25964, -29456, -30433, -30533, -30017, 
    -30629, -27059, -28326, -23989, -19889, -17384, -13145, -9331, -6451, 
    -2162, 2958, 8722, 12248, 15662, 19394, 23907, 25116, 26896, 28290, 
    29526, 30220, 30975, 30182, 30023, 25712, 24645, 21398, 18321, 13036, 
    8707, 5296, 291, -3247, -8631, -11535, -15199, -18927, -23272, -24232, 
    -27291, -30629, -30045, -31386, -31343, -30883, -27492, -27201, -24652, 
    -22516, -18576, -14716, -9825, -5398, -1179, 2849, 6175, 12015, 16525, 
    19418, 21107, 24639, 28043, 27260, 30744, 30772, 30326, 29286, 27357, 
    27380, 22671, 21096, 18359, 13819, 12033, 6620, 2705, -1988, -8381, 
    -10997, -13292, -18192, -21547, -26097, -28415, -27333, -29521, -31736, 
    -30381, -30389, -28623, -26927, -24416, -21533, -19382, -13854, -10912, 
    -5517, -2418, 3465, 6298, 10675, 16393, 18935, 21683, 24445, 28622, 
    27992, 29593, 30283, 31400, 28731, 29058, 27240, 24852, 21964, 17672, 
    13421, 10169, 5983, 3485, -1486, -6035, -10661, -15582, -18127, -20302, 
    -22866, -26796, -29476, -30033, -31650, -30656, -28569, -29578, -27619, 
    -26247, -21954, -17784, -14901, -11753, -7745, -3114, 338, 5785, 9867, 
    13017, 17913, 22396, 23837, 27765, 28275, 29535, 31028, 29918, 29676, 
    29084, 28547, 25038, 22898, 18036, 14576, 10719, 6536, 2840, -2492, 
    -4939, -9733, -12910, -17672, -21125, -24158, -26358, -28394, -29872, 
    -31536, -31855, -30097, -29172, -27546, -25271, -23378, -18377, -14781, 
    -11826, -7136, -2890, 1487, 5981, 9330, 13283, 17861, 19417, 25548, 
    27283, 29625, 29660, 29948, 30954, 30920, 28308, 27752, 24838, 23579, 
    19514, 15134, 11418, 7089, 1789, -1417, -5327, -9576, -12698, -18238, 
    -21657, -24522, -26612, -29091, -28874, -31064, -30109, -30009, -29834, 
    -27444, -24127, -22093, -20294, -16524, -12194, -8075, -2835, 804, 6274, 
    9642, 13244, 17068, 21646, 23432, 25793, 29098, 30713, 30149, 29935, 
    30918, 29361, 28424, 24821, 23085, 19651, 16661, 13190, 8997, 3808, -709, 
    -6317, -10248, -13484, -16118, -20991, -22799, -25845, -28547, -29427, 
    -30589, -30433, -30394, -28432, -27500, -25485, -23395, -19168, -16090, 
    -11403, -6968, -3116, -527, 4776, 8672, 12658, 18926, 20773, 22696, 
    25957, 28111, 28982, 30528, 30082, 29308, 31009, 27476, 24955, 21905, 
    20012, 16953, 11380, 7006, 4341, -257, -4501, -9448, -12987, -16717, 
    -19713, -24476, -26767, -27535, -28264, -29094, -30487, -30344, -28948, 
    -28757, -26992, -23289, -19347, -14909, -13561, -8437, -4970, -245, 4354, 
    7224, 13468, 16458, 21129, 22725, 25700, 27182, 29113, 30466, 30225, 
    31862, 29796, 28127, 26516, 23491, 20534, 15729, 11714, 8745, 5091, -982, 
    -4674, -9729, -12762, -18229, -20433, -23146, -25129, -27390, -28169, 
    -30452, -30104, -30020, -28422, -27184, -26409, -21774, -19355, -17387, 
    -11619, -10911, -3462, -1746, 4567, 6452, 12001, 15248, 18495, 22751, 
    26412, 27933, 29262, 30145, 29614, 29655, 30947, 29033, 25705, 23618, 
    21188, 17851, 12778, 9075, 6446, 855, -3844, -8700, -11687, -17126, 
    -19092, -23269, -24110, -29214, -30728, -30711, -29632, -31303, -30619, 
    -29656, -27249, -24963, -19222, -17210, -13878, -8249, -5991, -1872, 
    2831, 8664, 12028, 15020, 19251, 23149, 25137, 28813, 29062, 30385, 
    32238, 30237, 29594, 28497, 26262, 22632, 21202, 18577, 13263, 8608, 
    5238, 1307, -2948, -9164, -11614, -16110, -18115, -22603, -23902, -27711, 
    -29580, -31132, -30707, -31155, -29064, -27630, -27414, -24338, -20534, 
    -17208, -14672, -9349, -6581, -534, 2884, 5972, 12094, 16066, 18223, 
    22337, 25698, 26126, 29324, 30043, 31248, 30030, 28488, 28199, 28216, 
    25513, 21682, 17500, 14828, 10401, 5631, 1234, -3491, -6394, -11797, 
    -15049, -18686, -22333, -25420, -26916, -29411, -30352, -29741, -31018, 
    -29424, -29621, -27727, -25117, -21137, -18582, -14054, -9641, -5374, 
    -3072, 1374, 5400, 9842, 15412, 18810, 21005, 26024, 26270, 29330, 30705, 
    31731, 30899, 29922, 30582, 27866, 23972, 21938, 18359, 14767, 10290, 
    6208, 772, -788, -7027, -9686, -15994, -17405, -22132, -24744, -27233, 
    -28499, -30612, -29383, -31154, -29654, -28093, -27375, -24549, -21970, 
    -18392, -14717, -11661, -7205, -1718, 1171, 6849, 11681, 14185, 17613, 
    21927, 24416, 26364, 29457, 31179, 30271, 31018, 29128, 28008, 26954, 
    24717, 23070, 18691, 15681, 12059, 5994, 3064, -1014, -7586, -9961, 
    -15099, -18942, -21554, -25559, -26585, -28976, -30881, -31038, -29352, 
    -29745, -29018, -27589, -25680, -22757, -19208, -15460, -11134, -7075, 
    -2250, 890, 5840, 10887, 14788, 19718, 21545, 25331, 27460, 29432, 31212, 
    30929, 30765, 30512, 28338, 27761, 26682, 21363, 20332, 15233, 12906, 
    8051, 1944, 124, -6571, -10724, -14435, -18134, -21885, -24869, -27853, 
    -28121, -30188, -31755, -29845, -30321, -29447, -28049, -26359, -23987, 
    -17853, -16826, -12680, -9152, -2520, 1383, 5502, 9892, 13665, 16522, 
    20491, 23305, 27796, 29983, 28894, 29651, 32313, 30361, 29502, 27715, 
    24997, 22580, 20043, 16787, 11809, 8990, 2175, -630, -5343, -9618, 
    -14881, -17491, -20737, -24460, -27401, -29574, -29484, -31302, -31316, 
    -29755, -28612, -27667, -24246, -23556, -19911, -15560, -11044, -7374, 
    -2596, 124, 4743, 11023, 13060, 17532, 21964, 23319, 27259, 28181, 29231, 
    31226, 29023, 32096, 28566, 29070, 26126, 22725, 19035, 16246, 13465, 
    7428, 4222, -1507, -3676, -8493, -13369, -16096, -20709, -23415, -25429, 
    -27850, -30109, -30058, -30973, -29580, -29800, -27775, -24280, -23620, 
    -19717, -17052, -11656, -7357, -3714, 631, 5363, 8670, 12819, 17507, 
    19890, 23740, 27462, 27841, 30873, 30788, 31264, 29953, 28354, 28654, 
    25588, 23298, 20387, 15613, 12351, 8076, 4082, 862, -3578, -8831, -12284, 
    -16433, -19115, -24713, -25182, -26344, -30798, -31204, -31017, -30631, 
    -31034, -28053, -25242, -24318, -19730, -17142, -12827, -7988, -3817, 
    -1913, 3150, 8199, 11440, 17552, 19664, 24051, 27430, 28057, 29818, 
    31732, 31510, 31048, 30008, 28510, 26017, 24687, 22077, 16621, 13190, 
    7834, 4290, 1661, -3856, -7668, -13797, -16179, -19562, -22891, -26789, 
    -26705, -31018, -29870, -32012, -29698, -29861, -28754, -26228, -23825, 
    -19274, -17503, -13700, -8750, -3324, -541, 3748, 9377, 12476, 16582, 
    19507, 24321, 26616, 26797, 28486, 30133, 31137, 30305, 28932, 28566, 
    25566, 22978, 21183, 17782, 12095, 8638, 5020, 987, -4911, -9530, -12754, 
    -16027, -18758, -23287, -25500, -28380, -30873, -31872, -30623, -30255, 
    -28622, -27596, -25855, -24711, -21267, -18114, -12936, -9766, -5534, 
    368, 3041, 8768, 10982, 15871, 18568, 24191, 25443, 27914, 28754, 29756, 
    31751, 31545, 29672, 28526, 27232, 23740, 21492, 18710, 14120, 10353, 
    4387, 857, -4281, -7794, -11415, -14376, -19072, -22876, -25926, -26723, 
    -29590, -30188, -31444, -30367, -30490, -28792, -27764, -23291, -19996, 
    -18073, -13767, -8456, -5852, -1578, 4010, 7446, 10627, 15381, 20633, 
    21365, 25386, 26269, 28378, 29381, 29930, 31172, 29255, 29296, 26280, 
    24262, 21181, 18135, 13427, 9038, 6059, 1787, -2399, -7305, -11347, 
    -16140, -18245, -22727, -25705, -29077, -28349, -30526, -30155, -30495, 
    -30156, -27309, -27190, -24743, -20483, -18780, -13933, -10255, -4851, 
    -1750, 1977, 8539, 11115, 15402, 17941, 23228, 24679, 27366, 28598, 
    31012, 30887, 30499, 31084, 28064, 26365, 24422, 21410, 17247, 13758, 
    10259, 6950, 795, -3009, -6701, -11673, -14798, -19051, -21469, -24884, 
    -26633, -27770, -30711, -30215, -32103, -30279, -30532, -27159, -25656, 
    -21386, -19855, -13644, -10694, -6236, -3348, 2420, 6471, 10698, 15794, 
    19178, 22994, 23248, 27633, 27672, 30126, 30588, 30141, 31191, 28469, 
    25995, 23500, 20796, 18698, 13463, 10823, 7734, 2529, -2384, -6468, 
    -11645, -15773, -18021, -20933, -24154, -27034, -27852, -29716, -30880, 
    -30885, -29264, -29884, -26024, -24279, -23693, -19431, -14282, -10987, 
    -7541, -1661, 3317, 4918, 10142, 12767, 18718, 22006, 23267, 27253, 
    29432, 28730, 30387, 31644, 31173, 30830, 27856, 24247, 21079, 17304, 
    15280, 11116, 7339, 2701, -2387, -5835, -11802, -13635, -18021, -22565, 
    -25501, -27207, -28377, -29416, -29315, -31883, -30900, -29304, -26856, 
    -25431, -22369, -18811, -15649, -10787, -6861, -1844, 2256, 5084, 10366, 
    14638, 17816, 20464, 23409, 26953, 28076, 30467, 31770, 30898, 31228, 
    29678, 28175, 24834, 22590, 19459, 16214, 11426, 8604, 4081, -668, -5967, 
    -9744, -12560, -16013, -20403, -23624, -25562, -29800, -30984, -30952, 
    -30089, -29217, -29488, -27906, -26445, -21833, -19848, -17593, -11161, 
    -8117, -4148, 1145, 5180, 9609, 12384, 16202, 21268, 24268, 26261, 29360, 
    29394, 30589, 30474, 30475, 28284, 27012, 25850, 21159, 19248, 16356, 
    13586, 7917, 4785, -793, -3947, -8095, -12280, -16601, -19846, -23104, 
    -26888, -28810, -29844, -29277, -30419, -30774, -30134, -27139, -24998, 
    -24711, -20848, -16298, -12180, -9311, -3238, 680, 5226, 9820, 13856, 
    16754, 19761, 23573, 25169, 28583, 29372, 30266, 30106, 30671, 29379, 
    28335, 25144, 23987, 18844, 15563, 12439, 7674, 3573, -1481, -4721, 
    -9305, -13960, -16872, -19961, -23031, -26373, -27964, -28574, -30748, 
    -31237, -30764, -28767, -29205, -27409, -23002, -20757, -16581, -11047, 
    -6836, -3530, 204, 3617, 8957, 13354, 18052, 20207, 22578, 25286, 28874, 
    29925, 31180, 30286, 29730, 29280, 27955, 25817, 22271, 19207, 17414, 
    13992, 8826, 4667, 72, -4385, -9034, -12955, -17030, -19597, -23487, 
    -25191, -28326, -30900, -31653, -29741, -30430, -29768, -27617, -26348, 
    -22799, -19936, -17500, -14276, -8028, -3957, -1039, 2906, 8358, 11276, 
    16158, 20691, 22255, 24705, 27907, 29111, 29275, 29554, 30302, 29025, 
    28160, 26191, 23585, 21990, 17142, 12312, 8771, 4589, 505, -5038, -7473, 
    -11486, -15928, -20114, -22795, -25206, -28424, -28361, -30433, -31732, 
    -29714, -28638, -28260, -27581, -22822, -19466, -15905, -13446, -9219, 
    -6491, -1125, 3423, 7954, 11876, 15611, 20832, 22884, 25967, 27458, 
    29805, 31694, 30997, 30370, 29456, 28581, 26835, 23540, 19291, 18232, 
    14498, 8467, 5711, 1521, -2937, -7590, -10442, -14898, -20797, -23025, 
    -24156, -27562, -30250, -28799, -30765, -32019, -29779, -28652, -26719, 
    -24548, -20962, -18281, -13915, -11222, -5759, -967, 2291, 6826, 10828, 
    14702, 19318, 21210, 26057, 26914, 29918, 29157, 30806, 30865, 29728, 
    28197, 27330, 23590, 21783, 17435, 14629, 9365, 4064, 1237, -2387, -6043, 
    -11340, -16205, -18671, -20455, -24937, -27699, -27937, -29488, -32481, 
    -30057, -29764, -28802, -27222, -25337, -21030, -20015, -15427, -10013, 
    -6329, -609, 3554, 7179, 11469, 15488, 18727, 20729, 25353, 26022, 27703, 
    30046, 31572, 31116, 29205, 28816, 26503, 23086, 22236, 18438, 13900, 
    9821, 7767, 2511, -962, -5998, -11050, -14226, -18509, -21764, -23977, 
    -28028, -27722, -30597, -30855, -31038, -30272, -28951, -27817, -25639, 
    -21747, -18192, -14589, -9290, -7458, -1804, 654, 6148, 9424, 13932, 
    18172, 22038, 24410, 27152, 28517, 29872, 31809, 29668, 30805, 28351, 
    27935, 24468, 20730, 19811, 14972, 12721, 6357, 1353, -2432, -5144, 
    -10575, -14329, -18039, -21852, -23443, -25872, -29733, -30108, -29619, 
    -29866, -30106, -29734, -25958, -25033, -22219, -19066, -15610, -12141, 
    -7742, -3341, 3110, 6569, 9836, 12837, 17163, 22430, 24166, 27367, 27765, 
    28849, 30517, 32355, 30280, 29151, 25608, 24333, 22181, 19921, 15870, 
    11211, 5737, 4021, -2951, -7514, -8789, -15298, -17008, -21008, -22523, 
    -25825, -28714, -30933, -29182, -31413, -29378, -28956, -27562, -24583, 
    -22264, -20709, -14305, -11246, -6387, -4594, 509, 5875, 9088, 12937, 
    17006, 22771, 23707, 25525, 28345, 31470, 29322, 30777, 30255, 30309, 
    25951, 25434, 23667, 19462, 16965, 12834, 8201, 2789, -1082, -6651, 
    -10243, -13638, -16954, -21198, -22831, -26097, -26926, -28926, -31537, 
    -32473, -30274, -30488, -28134, -25786, -22703, -19526, -15633, -12612, 
    -8840, -3759, 1825, 5897, 9087, 13219, 15905, 20295, 23386, 26984, 28459, 
    30074, 30245, 30784, 28514, 29189, 26663, 24837, 24582, 19557, 15844, 
    12627, 7539, 3724, -496, -4244, -10161, -14185, -17632, -20879, -24558, 
    -24732, -28148, -30538, -32054, -31395, -30549, -28418, -27367, -26126, 
    -22236, -21086, -16751, -13146, -7638, -4340, 385, 4670, 9692, 12702, 
    17178, 20319, 23550, 26425, 28363, 28730, 31049, 29964, 31084, 28309, 
    28084, 26879, 24644, 21380, 15267, 12407, 6960, 5380, 418, -3970, -9057, 
    -13994, -17773, -20033, -25063, -26347, -28217, -30153, -31173, -30440, 
    -31100, -30531, -28720, -26771, -22608, -20378, -17721, -13697, -8444, 
    -4606, 552, 3320, 8428, 13658, 17538, 20317, 22807, 25176, 26933, 29699, 
    29793, 29627, 29832, 28129, 26602, 26485, 23374, 21347, 15112, 14266, 
    9334, 4225, -963, -3892, -8409, -13925, -16351, -21785, -23773, -26018, 
    -27488, -30664, -31061, -30850, -30417, -29805, -27782, -27156, -24510, 
    -21415, -17216, -13152, -8007, -5076, -796, 2738, 9423, 12719, 14358, 
    18716, 21614, 26674, 27432, 29149, 28931, 30743, 30121, 31012, 28925, 
    25028, 24898, 21412, 17432, 13619, 8885, 3456, 1823, -4881, -8750, 
    -13223, -16272, -18970, -21749, -26697, -28194, -29536, -30795, -30337, 
    -29260, -28881, -28371, -27813, -23986, -20392, -16421, -12725, -9482, 
    -4772, -208, 3644, 6607, 10894, 14345, 19352, 21513, 23666, 27285, 27916, 
    31131, 31346, 29379, 29148, 28959, 26277, 22846, 21362, 17415, 13118, 
    9609, 3848, 2163, -2040, -8282, -12366, -16885, -20041, -21730, -26011, 
    -26474, -28714, -29801, -30781, -29961, -30026, -27989, -25935, -24867, 
    -22374, -19588, -12980, -9138, -5775, -1311, 4253, 7225, 11470, 14567, 
    19891, 21916, 23789, 26751, 30115, 28782, 31234, 30176, 28935, 28911, 
    27969, 23626, 22290, 17195, 14722, 10171, 5767, 2434, -3831, -7748, 
    -10537, -14764, -19133, -22828, -24946, -26276, -29417, -29853, -30872, 
    -32347, -29457, -29052, -26952, -24490, -21540, -17551, -15200, -10725, 
    -4641, -1746, 1306, 6283, 11588, 15997, 19186, 22255, 24140, 27442, 
    29619, 31886, 30335, 31429, 30152, 28778, 26507, 24514, 21826, 19720, 
    15139, 9676, 6825, 2539, -3068, -8076, -11404, -14675, -17099, -21551, 
    -25327, -26518, -29417, -29775, -28944, -30138, -29675, -29217, -27446, 
    -25146, -22731, -18380, -13542, -11191, -5687, -1949, 2299, 7162, 10805, 
    15218, 18329, 21691, 24233, 26436, 29083, 31331, 30493, 30796, 29930, 
    28991, 26989, 26243, 22455, 18272, 14420, 11042, 6808, 3505, -2852, 
    -6521, -9909, -13841, -17807, -21078, -25863, -28185, -28528, -30333, 
    -30187, -31161, -30870, -29678, -27727, -24665, -20723, -18285, -16827, 
    -10196, -7552, -2781, 2242, 6736, 11434, 13120, 19266, 22223, 24849, 
    27416, 29333, 29702, 30923, 30445, 30110, 28658, 27499, 25667, 21891, 
    18520, 14330, 12196, 8242, 2826, -2153, -4973, -10664, -15825, -19067, 
    -21591, -24499, -28290, -28795, -29917, -31031, -31397, -30605, -28421, 
    -27356, -24966, -22748, -17680, -14447, -12354, -7742, -1664, 2677, 7248, 
    10585, 13391, 17098, 21600, 24474, 27976, 27976, 30779, 29009, 30705, 
    28573, 29165, 28162, 25431, 24320, 19295, 14291, 10410, 8692, 2916, 
    -1328, -7095, -9893, -13821, -17658, -22745, -23198, -26008, -27348, 
    -30420, -31201, -30330, -31763, -29493, -28981, -23581, -20960, -18329, 
    -16624, -12453, -7652, -4799, 1063, 6293, 9245, 14705, 17174, 19353, 
    24968, 25907, 27261, 30510, 30350, 30986, 31470, 29518, 28073, 25675, 
    22010, 20058, 14622, 11962, 8128, 3533, -342, -6209, -8963, -13295, 
    -18730, -20797, -23492, -27327, -27280, -29987, -30745, -29303, -29594, 
    -29451, -29017, -27087, -23702, -20943, -17405, -12261, -8357, -4844, 
    1065, 3822, 9182, 12135, 18629, 20384, 23127, 26921, 27829, 30815, 31102, 
    30223, 29968, 30912, 27555, 24947, 23092, 20140, 17334, 12187, 8029, 
    3433, -1359, -4791, -8960, -12338, -16531, -19834, -24465, -26876, 
    -27598, -29864, -31400, -30330, -30342, -29551, -26320, -26108, -23118, 
    -19420, -18389, -12557, -6897, -3802, -982, 2821, 9386, 13613, 16897, 
    20597, 23161, 26620, 27818, 29573, 30922, 30718, 30938, 29147, 27989, 
    24545, 24416, 19419, 16746, 13876, 9996, 3483, -181, -3330, -9646, 
    -11689, -16440, -20154, -23157, -27165, -27285, -28140, -30696, -31546, 
    -29543, -30925, -27446, -25259, -23503, -18847, -16030, -13428, -8592, 
    -5294, -940, 3690, 7840, 13185, 15462, 19234, 23390, 26985, 29263, 29569, 
    29889, 31770, 30799, 29904, 27278, 26511, 22810, 20462, 18737, 14120, 
    10011, 5405, 2442, -3295, -6949, -11610, -16676, -18792, -23244, -27209, 
    -27890, -29486, -30134, -30882, -31641, -30268, -29104, -24952, -23489, 
    -20977, -18550, -13078, -8743, -5367, -1354, 3931, 8646, 12320, 15705, 
    19080, 23872, 25142, 26508, 29461, 30772, 30608, 31616, 30458, 28422, 
    27288, 23893, 20463, 16781, 13985, 9669, 4199, 2556, -2801, -6500, 
    -11214, -15745, -18318, -22804, -25244, -26891, -28221, -30250, -30249, 
    -29251, -31543, -28261, -25107, -23988, -19903, -16727, -13006, -9798, 
    -7120, -1181, 3235, 7282, 11621, 16026, 20337, 21853, 24982, 27167, 
    27865, 31081, 32552, 29536, 30097, 28184, 26398, 23216, 20179, 18018, 
    14091, 9470, 7276, 137, -2494, -8481, -10195, -16502, -18621, -22025, 
    -23883, -27107, -28744, -30066, -30474, -29567, -29008, -28886, -27371, 
    -24960, -21539, -17333, -15837, -9875, -4717, -1549, 4134, 6459, 11744, 
    14343, 19857, 22285, 24974, 27916, 28887, 30189, 31520, 29893, 30308, 
    28568, 26905, 25759, 22689, 18300, 13593, 9368, 6494, 1845, -2192, -6591, 
    -11079, -15132, -18898, -21663, -26022, -27129, -29559, -28938, -30627, 
    -30720, -31571, -29710, -28115, -24603, -20822, -16826, -13960, -9226, 
    -6750, -2267, 2505, 6250, 9956, 14002, 17644, 22607, 24915, 26706, 29703, 
    30143, 30893, 30800, 30606, 28417, 27580, 26091, 21907, 19524, 14505, 
    10798, 6040, 3842, -1899, -6912, -10265, -13967, -18186, -22000, -25418, 
    -27821, -29139, -30868, -29754, -29723, -31244, -29999, -25538, -24867, 
    -22173, -18285, -15579, -11393, -5680, -2741, 2820, 5370, 9796, 13648, 
    19011, 22287, 24426, 26742, 29010, 30148, 30823, 29520, 29709, 28074, 
    26264, 24967, 21744, 19250, 15839, 12373, 9022, 3290, -1364, -6458, 
    -9016, -13370, -18322, -20335, -24952, -27612, -30363, -29844, -31069, 
    -30888, -30402, -29956, -27230, -25799, -23505, -19652, -14854, -11214, 
    -6056, -3328, 1819, 5875, 10842, 14098, 18730, 20229, 24856, 26334, 
    29158, 30285, 30619, 32263, 30093, 29726, 26623, 26002, 23665, 19296, 
    14998, 10937, 7466, 3531, -137, -5239, -11305, -13867, -17667, -22573, 
    -24279, -26080, -27902, -28719, -31049, -29486, -30648, -29663, -27149, 
    -26178, -24047, -18064, -15048, -10551, -8539, -3344, 864, 3759, 9626, 
    13079, 15812, 19468, 22916, 27737, 28099, 28916, 30646, 30452, 30429, 
    29456, 28866, 26030, 23494, 18268, 14543, 11839, 8752, 3226, -1975, 
    -3278, -8567, -12902, -16996, -20308, -23530, -27991, -27242, -29414, 
    -30430, -30856, -31896, -28535, -27768, -26613, -22919, -20427, -17142, 
    -13096, -7987, -3404, 297, 4337, 7850, 13079, 18076, 21650, 23268, 26041, 
    28330, 31268, 29852, 30936, 29177, 28242, 27760, 26350, 23258, 19171, 
    16802, 11526, 9089, 4447, -317, -3937, -7668, -11810, -16126, -20878, 
    -21647, -26472, -27214, -29437, -32049, -31135, -29979, -31071, -27735, 
    -25330, -24054, -19565, -16725, -13864, -7603, -4369, -835, 4097, 8459, 
    13152, 17078, 19098, 23413, 26741, 27850, 30307, 30586, 31269, 31581, 
    28882, 27657, 26009, 23139, 20994, 17992, 12672, 9247, 4742, 774, -4115, 
    -6925, -13546, -16887, -19588, -24937, -25523, -28320, -28624, -29486, 
    -31523, -30298, -29764, -29441, -26117, -24081, -19387, -16918, -14420, 
    -8290, -4859, -1692, 3178, 9269, 11930, 16989, 21369, 23371, 25900, 
    28135, 29904, 29302, 31460, 30931, 30491, 27850, 26243, 22637, 19497, 
    17408, 13563, 8459, 4258, 185, -2437, -7538, -13150, -16849, -19072, 
    -23061, -26095, -27905, -28553, -31149, -31640, -30875, -29327, -29602, 
    -27309, -24044, -21710, -16509, -13316, -10151, -5040, -878, 3722, 7791, 
    12042, 16300, 19122, 23198, 24786, 26086, 28626, 30142, 31605, 30118, 
    30257, 28857, 26671, 25135, 21140, 18345, 14508, 9463, 6535, 1148, -2094, 
    -8075, -11995, -15198, -18042, -21879, -26254, -27493, -28609, -30445, 
    -29212, -29182, -30580, -27799, -26822, -24093, -21309, -18021, -14540, 
    -10595, -5109, -134, 1960, 7497, 12442, 16311, 19433, 21973, 24613, 
    28785, 28316, 30784, 31015, 31651, 28637, 28494, 26821, 24507, 21543, 
    16882, 14001, 9473, 5223, 508, -2505, -7170, -11145, -15211, -19953, 
    -20424, -25725, -27009, -28314, -28905, -31896, -29490, -30380, -29691, 
    -27662, -22566, -22855, -18773, -13079, -10693, -6189, -2693, 1140, 8052, 
    11880, 13535, 18415, 22122, 24676, 26981, 30526, 29205, 30692, 31030, 
    30155, 29105, 27188, 24245, 22323, 19323, 14160, 12034, 5304, 2776, 
    -3134, -6740, -11053, -15552, -16906, -21380, -25088, -27248, -30184, 
    -30638, -30729, -31248, -31734, -29312, -28367, -25258, -21403, -17954, 
    -14056, -12312, -7812, -2387, 2632, 6738, 9939, 14964, 18047, 21608, 
    23881, 28321, 28581, 29948, 29544, 29110, 30109, 28781, 25900, 25040, 
    22176, 18350, 15941, 11189, 6878, 2588, -1946, -5951, -9767, -13728, 
    -18707, -22633, -25450, -27011, -29431, -29501, -32351, -29611, -31107, 
    -30752, -27561, -24096, -22236, -18393, -15406, -11846, -5908, -2402, 
    409, 7140, 11494, 13975, 17276, 21157, 25671, 25976, 30235, 30477, 31732, 
    30341, 31915, 27621, 28520, 25454, 21086, 17260, 15810, 12078, 7921, 
    1663, -2139, -5396, -11376, -15838, -16366, -20959, -22797, -26537, 
    -27512, -29797, -29553, -30068, -31454, -29487, -27020, -26818, -22332, 
    -19054, -16284, -11918, -8758, -3409, 2254, 5995, 9295, 14324, 18152, 
    21314, 23056, 27001, 27397, 30361, 30233, 30828, 30882, 29637, 28190, 
    26013, 22108, 18763, 15534, 12197, 8483, 3902, -1873, -5922, -9636, 
    -13797, -17964, -22032, -24181, -25629, -28636, -30531, -30574, -30502, 
    -30490, -29191, -27484, -26895, -21448, -19707, -16281, -12201, -6806, 
    -1929, -34, 6743, 8819, 14812, 17905, 18987, 23942, 25827, 29475, 30249, 
    30724, 31147, 30582, 28617, 28065, 26970, 22926, 19083, 15947, 13243, 
    6641, 4162, -5, -6008, -9045, -13554, -17008, -21760, -23598, -26103, 
    -29013, -29578, -30622, -30964, -30806, -29882, -28807, -26413, -22058, 
    -20237, -15096, -12365, -9007, -4694, -698, 5390, 9884, 14816, 17991, 
    21005, 23519, 25828, 28231, 30386, 30275, 29274, 29561, 30432, 26326, 
    25585, 22504, 21049, 17994, 13063, 7560, 5709, -406, -3512, -9458, 
    -13276, -15662, -21151, -23052, -25057, -29875, -30298, -30491, -32253, 
    -31065, -30145, -28682, -26402, -21989, -20459, -18529, -13600, -7777, 
    -4640, 877, 5046, 9160, 13513, 17128, 20272, 22797, 25427, 28227, 28599, 
    30550, 32432, 30881, 30145, 27919, 26536, 23335, 19467, 15518, 12642, 
    8745, 4132, 752, -3723, -8681, -13105, -15449, -20286, -22995, -26066, 
    -29653, -29186, -30413, -31105, -29311, -29852, -29593, -25428, -25022, 
    -20392, -15827, -12816, -8555, -4058, -14, 2757, 8005, 12515, 15512, 
    20008, 21391, 27047, 28187, 29504, 31075, 29590, 29820, 29469, 28589, 
    24610, 23513, 20994, 16718, 12909, 8150, 5769, 1981, -4602, -9438, 
    -11815, -14259, -18611, -22991, -25644, -28260, -29273, -30231, -31416, 
    -30676, -29486, -28794, -26422, -22852, -21048, -17726, -14836, -9321, 
    -5130, -442, 3058, 8187, 12172, 16580, 18641, 23436, 24177, 27160, 27933, 
    29806, 31506, 30206, 30394, 29535, 25809, 23841, 20771, 18467, 12990, 
    9817, 4816, 391, -1916, -7408, -11703, -15507, -19585, -22846, -23480, 
    -26031, -28771, -30049, -30675, -30296, -29938, -28189, -28500, -24159, 
    -21791, -17285, -13990, -9751, -4897, -698, 3848, 7084, 11289, 16653, 
    19488, 21621, 26848, 28227, 28804, 30967, 32550, 29214, 30291, 28268, 
    25179, 24763, 21327, 17090, 13802, 9643, 4664, 2975, -2658, -8852, 
    -12327, -16387, -18349, -22296, -25407, -27075, -29602, -29424, -32167, 
    -29755, -30848, -29149, -26971, -23917, -22095, -17250, -15036, -11136, 
    -6228, -2032, 1196, 7975, 12185, 15440, 20500, 21560, 24412, 26187, 
    27648, 31053, 32258, 30775, 30126, 28378, 26949, 24725, 19902, 18625, 
    13391, 11714, 5705, 2388, -2003, -6033, -10547, -14120, -19024, -21167, 
    -23519, -27518, -28950, -28996, -30435, -30688, -29445, -29767, -27497, 
    -25682, -21822, -19050, -15732, -10971, -5961, -2930, 1442, 6503, 9695, 
    14432, 17124, 22925, 23638, 27807, 27565, 29580, 31183, 31341, 30519, 
    29435, 27217, 23903, 22493, 17537, 15396, 11148, 6269, 2758, -1577, 
    -7489, -10774, -14624, -19429, -21973, -25377, -27586, -28785, -30651, 
    -30278, -30831, -31518, -28431, -27671, -25467, -22006, -18101, -15127, 
    -11618, -6856, -1720, 1725, 5818, 8891, 14783, 18308, 21455, 24124, 
    26870, 28494, 31599, 32043, 30393, 31222, 29952, 27285, 25494, 22421, 
    19615, 15638, 11402, 6930, 2295, -2942, -4678, -8503, -14456, -17714, 
    -21345, -25381, -26657, -28372, -28456, -31252, -32192, -31787, -29816, 
    -28228, -25278, -22220, -19037, -16531, -11966, -6705, -1585, 1096, 4022, 
    11163, 14709, 19229, 22157, 22395, 25383, 27649, 30275, 30695, 30770, 
    30100, 29919, 28977, 24856, 23135, 17775, 15431, 11975, 8536, 2576, 
    -1578, -5185, -9296, -14342, -17484, -21366, -23284, -26599, -28929, 
    -29241, -30127, -30285, -31680, -29986, -27275, -23809, -22328, -20332, 
    -15406, -11258, -7370, -4421, -477, 6385, 9566, 12249, 16329, 20924, 
    23265, 25157, 27242, 29801, 31880, 30718, 29395, 28914, 27568, 25380, 
    23583, 19805, 16932, 13089, 7787, 1829, -760, -4224, -9401, -11821, 
    -15957, -20015, -23748, -27799, -27122, -30887, -31654, -31075, -30393, 
    -29205, -28582, -27051, -22763, -20784, -16913, -13372, -8752, -3235, 
    249, 5994, 8942, 13346, 17936, 20633, 23514, 26660, 28140, 30905, 29503, 
    31020, 29855, 27645, 29456, 24708, 22535, 19309, 16038, 12129, 9808, 
    3268, -681, -5212, -9882, -11845, -17845, -21551, -22786, -25692, -28464, 
    -30279, -30601, -31451, -31979, -29666, -27065, -26349, -23366, -18700, 
    -16999, -12176, -9078, -4156, 59, 4712, 8623, 14189, 17514, 19566, 22300, 
    25453, 28823, 29449, 31117, 31907, 32152, 30938, 26626, 25758, 24377, 
    18613, 16199, 13184, 9175, 5449, 281, -3897, -7928, -12621, -16703, 
    -20156, -21899, -25258, -28174, -27846, -31251, -31305, -31544, -29821, 
    -27766, -25545, -22709, -21311, -17024, -12346, -7624, -4285, 376, 4519, 
    7970, 12234, 14992, 20718, 23280, 25636, 27782, 30131, 29452, 31442, 
    30023, 30814, 28897, 27794, 23026, 20089, 18401, 12792, 9293, 3810, -42, 
    -2135, -8063, -11362, -15615, -20983, -23264, -24909, -27500, -28689, 
    -30440, -30538, -31091, -28941, -28419, -27773, -23708, -21602, -17487, 
    -13730, -7916, -6891, 443, 4177, 7547, 12823, 16218, 19240, 22683, 25572, 
    27369, 28580, 29840, 31171, 30151, 29879, 27687, 26758, 24234, 20893, 
    16514, 12415, 8255, 5319, 1783, -2710, -8596, -12483, -15347, -20906, 
    -21516, -26137, -27196, -28669, -30230, -30447, -30569, -28237, -27754, 
    -26645, -24216, -20350, -18072, -13727, -9756, -6044, -314, 3199, 7855, 
    12017, 16418, 18547, 22128, 24539, 27413, 27929, 30468, 31593, 30740, 
    29254, 29257, 26751, 24655, 22755, 17408, 12919, 11447, 5705, 2381, 
    -2701, -7974, -10978, -14624, -18873, -23231, -24204, -27340, -28174, 
    -31642, -31694, -31080, -28602, -28447, -27057, -23614, -21434, -18190, 
    -13984, -11462, -4770, -2315, 3380, 7599, 11989, 16163, 18738, 23472, 
    24982, 28107, 27746, 29390, 31019, 30702, 29630, 27196, 25792, 25401, 
    21856, 17822, 16347, 10587, 7040, 1959, -2878, -5809, -11324, -14797, 
    -19004, -22193, -24580, -25661, -28882, -30820, -30841, -30791, -30783, 
    -28919, -27640, -24074, -21795, -19917, -14021, -10629, -6452, -2487, 
    4017, 7269, 10631, 13563, 18116, 21245, 26526, 28493, 27982, 31037, 
    31719, 30586, 29877, 28879, 28266, 23735, 21532, 19634, 13612, 10912, 
    7607, 2560, -2040, -6313, -9894, -13330, -18601, -21785, -24903, -26107, 
    -29073, -29263, -30953, -31060, -30199, -29209, -26984, -24535, -23266, 
    -17860, -15040, -11234, -6751, -3046, 523, 6429, 10151, 15389, 18143, 
    21791, 23367, 26432, 28559, 30872, 30041, 29123, 31015, 28914, 27768, 
    23714, 23119, 17413, 16402, 11191, 6828, 3897, -1551, -6700, -10925, 
    -15262, -18037, -20948, -24609, -26479, -29146, -30976, -31339, -31377, 
    -29740, -29553, -28420, -24878, -21564, -18619, -14501, -11767, -7373, 
    -3275, 1995, 4406, 9610, 12737, 18152, 21113, 24518, 25827, 28481, 28700, 
    31304, 30964, 29965, 30742, 26359, 24973, 22146, 18558, 16670, 12436, 
    7779, 2571, -2599, -5471, -9911, -14058, -17516, -22005, -25343, -26028, 
    -27882, -30355, -29383, -30618, -29732, -29466, -27813, -24749, -21033, 
    -18014, -16737, -13305, -7005, -3471, -280, 6312, 8646, 12564, 17385, 
    21112, 23036, 25908, 28336, 29838, 31163, 30588, 30324, 28843, 28086, 
    24622, 23468, 20139, 15638, 12510, 7539, 2468, -1987, -5387, -8609, 
    -11824, -16279, -19517, -24088, -25729, -28951, -29729, -30713, -30746, 
    -30054, -29248, -27077, -26770, -24605, -19575, -14903, -12496, -8285, 
    -3536, 1233, 5265, 10703, 14322, 16503, 21997, 23054, 25543, 28430, 
    28309, 29544, 30738, 29313, 29346, 28123, 24482, 22877, 20308, 17293, 
    11916, 8450, 5242, -70, -5255, -7157, -12791, -16163, -18808, -24259, 
    -27122, -28419, -30167, -30629, -31255, -28832, -30023, -28762, -24686, 
    -22311, -20515, -16158, -12550, -9705, -3967, -177, 4938, 8288, 13309, 
    16715, 20068, 23593, 25143, 28370, 30359, 30467, 29241, 31461, 31273, 
    28657, 26192, 23224, 19444, 17550, 11313, 9440, 4204, -1418, -3859, 
    -8413, -13398, -15935, -19972, -22015, -25791, -28062, -30573, -31054, 
    -31904, -29425, -30380, -29165, -26961, -23024, -19535, -16822, -13324, 
    -9669, -5453, -162, 2752, 8564, 13259, 14493, 18592, 23237, 24189, 28122, 
    28904, 29732, 30632, 30711, 28686, 28968, 25805, 24759, 20842, 16223, 
    14390, 8532, 4916, -386, -4370, -9092, -12295, -17789, -19853, -22237, 
    -24775, -27738, -29155, -30727, -30079, -30378, -29347, -27498, -26465, 
    -24507, -21250, -16862, -13541, -9096, -5000, -1201, 3667, 7908, 13178, 
    15258, 20718, 22415, 26042, 26626, 29970, 31284, 32006, 30886, 29826, 
    28692, 27363, 22795, 21195, 18799, 12763, 8750, 4502, 1685, -3713, -7009, 
    -13076, -16810, -18416, -21914, -25132, -26045, -29334, -29507, -30314, 
    -31420, -29829, -27751, -27003, -22812, -19716, -19340, -13526, -8652, 
    -6205, -1826, 2421, 6807, 11186, 15478, 19953, 23215, 24779, 27701, 
    30043, 30021, 31740, 30720, 29138, 28618, 26800, 24293, 21963, 18303, 
    15074, 9937, 7386, 2157, -3788, -6816, -9968, -14271, -19763, -21253, 
    -24786, -27299, -28592, -31214, -30979, -30240, -28932, -27439, -27562, 
    -24100, -21309, -16732, -14508, -10397, -6651, -1905, 4116, 6784, 11759, 
    15378, 17368, 20973, 24582, 27969, 29878, 29137, 29911, 31694, 29323, 
    29060, 26487, 25104, 22775, 17466, 13428, 9795, 5576, 304, -1792, -6813, 
    -10977, -15842, -18091, -21648, -23655, -25657, -29221, -29456, -30882, 
    -31386, -30163, -28218, -26489, -25871, -21442, -18541, -14541, -10161, 
    -7196, -2562, 1591, 6821, 11105, 13664, 18877, 22558, 25607, 27629, 
    28380, 29739, 30209, 29868, 29885, 29691, 27892, 25596, 22100, 17402, 
    15405, 10288, 7041, 2033, -2414, -5677, -10955, -14768, -17161, -22216, 
    -25409, -26668, -30098, -28933, -32473, -30408, -28899, -29490, -28101, 
    -25864, -20658, -19160, -14629, -9875, -6182, -756, 884, 5135, 9272, 
    13447, 18437, 21430, 24907, 25187, 29604, 29713, 31625, 30514, 30718, 
    28891, 27649, 24410, 23291, 19365, 15361, 11875, 7236, 2683, -1354, 
    -7728, -9871, -14374, -17242, -20686, -24152, -26540, -28686, -30305, 
    -29990, -31510, -31378, -30277, -28386, -23694, -21752, -20628, -15601, 
    -10913, -7744, -3777, 1498, 6308, 10090, 14033, 17662, 20792, 24634, 
    27244, 29832, 29877, 29378, 31201, 31347, 30385, 28689, 25338, 22621, 
    20226, 15747, 11173, 8743, 2430, -449, -5358, -10181, -14144, -16106, 
    -20614, -24630, -26895, -29321, -29140, -29171, -30716, -31420, -27671, 
    -26481, -24895, -23501, -20894, -15491, -11853, -7274, -3425, 1468, 4591, 
    8994, 13939, 15844, 21289, 24249, 26711, 29427, 29917, 30899, 29637, 
    31593, 29952, 27553, 24286, 22119, 19098, 16875, 11705, 7369, 3674, 
    -1864, -4713, -10804, -13783, -18334, -19637, -24052, -26666, -28705, 
    -30897, -30557, -32555, -30406, -29416, -26892, -26032, -22652, -20058, 
    -15179, -12514, -8483, -3142, -10, 3664, 9486, 13387, 16930, 19843, 
    23845, 25237, 28673, 29689, 30534, 31040, 29841, 28867, 26503, 24888, 
    24425, 21544, 15884, 12814, 8874, 4073, -873, -5211, -7403, -11920, 
    -15901, -19618, -23567, -26160, -29045, -29478, -30725, -30306, -30505, 
    -30006, -26673, -27497, -22232, -19326, -16716, -12674, -9823, -4809, 
    -452, 2859, 8032, 14371, 16602, 19721, 25098, 24043, 26977, 30016, 30372, 
    31685, 30516, 29354, 27650, 26444, 23268, 19975, 16912, 11673, 8261, 
    4643, -465, -4798, -8721, -13069, -17870, -19750, -22702, -25755, -26466, 
    -29016, -29893, -31437, -30357, -30045, -28337, -25422, -22841, -20441, 
    -16347, -13208, -8927, -5776, -196, 2348, 9567, 12497, 16103, 20622, 
    21971, 25963, 29403, 29118, 31470, 31140, 31659, 29575, 28520, 24967, 
    24552, 20210, 17438, 14540, 9424, 3754, 759, -3776, -8673, -11775, 
    -16426, -17949, -24046, -25109, -27060, -29213, -30242, -31039, -30948, 
    -30830, -29947, -27383, -24163, -19783, -17415, -13820, -9442, -4102, 
    -1231, 1987, 7523, 11609, 16080, 19991, 22064, 25291, 27430, 28290, 
    30399, 30379, 31429, 29758, 28817, 25400, 24210, 20897, 19414, 14486, 
    9303, 6198, 2699, -3256, -7540, -12221, -15594, -18548, -22829, -24773, 
    -28493, -28676, -28928, -32406, -30306, -29427, -27354, -27805, -25004, 
    -22381, -18511, -15165, -10877, -4329, -684, 3597, 8081, 12707, 15847, 
    19631, 20800, 26338, 27806, 29286, 28911, 31392, 32194, 30110, 28937, 
    26143, 24433, 21605, 18535, 13337, 10711, 6495, 1283, -4124, -8359, 
    -11366, -15724, -19100, -22285, -24424, -27322, -28732, -31006, -29218, 
    -30356, -29748, -30507, -28513, -25775, -21435, -19592, -13656, -10594, 
    -6232, -344, 1063, 5348, 10135, 14041, 20217, 21805, 24553, 28463, 29307, 
    29533, 30446, 30520, 30146, 27948, 26430, 26091, 20722, 18271, 13959, 
    11365, 6714, 1063, -2576, -6050, -11769, -14035, -19057, -22277, -23510, 
    -28770, -27989, -29785, -30990, -30641, -28887, -27796, -28714, -25610, 
    -21064, -18864, -14277, -12105, -7644, -1119, 3018, 6568, 10589, 14663, 
    19162, 21784, 26032, 26966, 27142, 28709, 32259, 30010, 31440, 28913, 
    27360, 24558, 22568, 18177, 14040, 11855, 6584, 3979, -1717, -6151, 
    -9592, -15338, -19195, -22010, -24338, -27813, -29076, -30456, -30661, 
    -30322, -29185, -28608, -27103, -23884, -22636, -17938, -14710, -10550, 
    -5852, -3809, 2541, 6333, 8925, 15131, 17756, 22141, 23789, 26553, 28844, 
    30850, 30631, 30315, 30182, 28144, 26642, 24487, 20705, 19171, 14906, 
    11459, 6723, 3504, -2243, -7147, -10329, -14114, -17663, -21298, -23981, 
    -25755, -28370, -29465, -31026, -30639, -29414, -28631, -28335, -24140, 
    -23240, -17736, -15221, -11690, -7226, -2589, 2744, 4999, 10078, 15207, 
    18071, 20679, 24066, 26114, 27623, 30793, 31370, 29288, 28658, 29254, 
    26434, 26889, 23538, 20604, 16239, 11270, 7506, 3528, -1400, -6574, 
    -8068, -12044, -18159, -20364, -24156, -25889, -27556, -29400, -28836, 
    -30107, -30034, -28124, -28635, -26835, -22394, -20731, -15421, -10570, 
    -8212, -2309, 1061, 5244, 9717, 13814, 17458, 22242, 23582, 27198, 27989, 
    28819, 30003, 30451, 30718, 29497, 27113, 25444, 23034, 20664, 16166, 
    12927, 7439, 3749, -200, -5688, -9962, -12717, -17227, -20120, -24112, 
    -27721, -28240, -29067, -30553, -29911, -29243, -29286, -27128, -26489, 
    -21499, -20051, -15420, -11489, -9812, -3238, 249, 6178, 7427, 13109, 
    16148, 19713, 23194, 26926, 28574, 29642, 31784, 32526, 30916, 28970, 
    28309, 25640, 23229, 20246, 16677, 12985, 8821, 3990, 558, -4899, -8689, 
    -12927, -17293, -19078, -21760, -25557, -28928, -29604, -29640, -30047, 
    -29212, -28294, -27954, -24837, -23754, -20185, -17426, -13467, -9256, 
    -3765, 1432, 4769, 9712, 12356, 16599, 19244, 21682, 25952, 27792, 31177, 
    30386, 30100, 30374, 29574, 27542, 26525, 23539, 20465, 16895, 12341, 
    9314, 4165, -144, -3559, -9845, -11940, -16881, -20409, -23077, -27007, 
    -26426, -29434, -31053, -29873, -31145, -29175, -29248, -25051, -22913, 
    -21233, -18169, -11753, -9653, -5565, 511, 4538, 7226, 13008, 16541, 
    20280, 22605, 26243, 29021, 28385, 30811, 31323, 30800, 29647, 28054, 
    27198, 24917, 21640, 17531, 13518, 8593, 5680, 1417, -4152, -7312, 
    -11559, -16839, -20112, -22839, -25344, -29365, -29405, -31469, -31056, 
    -30842, -31001, -28188, -26430, -25553, -21134, -17296, -13408, -8724, 
    -5618, -323, 4336, 7893, 11587, 17042, 20382, 23215, 24464, 27803, 30247, 
    31012, 30401, 29924, 29728, 26746, 27026, 23844, 19845, 19007, 13575, 
    8636, 6537, 641, -3339, -7738, -12755, -15427, -18944, -22762, -24800, 
    -27504, -28710, -29183, -31311, -30273, -29137, -28430, -27376, -23303, 
    -20330, -18537, -14533, -9430, -6216, -1021, 2192, 7347, 11557, 16535, 
    19544, 22302, 24329, 27710, 27629, 30221, 32105, 30099, 30097, 28836, 
    27280, 23348, 22416, 17174, 14025, 9706, 5659, 2178, -2953, -6881, 
    -12797, -15504, -19323, -20981, -23624, -27624, -29060, -30580, -30265, 
    -32162, -28640, -28626, -26883, -23870, -23034, -17712, -14866, -9678, 
    -6020, -2877, 2550, 5520, 11379, 15985, 18219, 21728, 23193, 26570, 
    28715, 29020, 31055, 30828, 29753, 28968, 26494, 24081, 22152, 17946, 
    12760, 11608, 6722, 2028, -2008, -7273, -10648, -14752, -18802, -21451, 
    -24805, -27696, -29632, -29902, -30003, -29225, -30962, -28900, -26539, 
    -24232, -21470, -18440, -15419, -11976, -5210, -2367, 1641, 5265, 11499, 
    15807, 18707, 21645, 23421, 27474, 29814, 30891, 31372, 30556, 30736, 
    28805, 26966, 24645, 21563, 20384, 14955, 10634, 5985, 4146, -2829, 
    -7215, -10895, -13853, -17651, -20499, -25919, -26518, -28322, -30307, 
    -32185, -30814, -30824, -28107, -27158, -23202, -21436, -17265, -14630, 
    -10233, -7227, -1050, 3496, 6602, 9209, 14241, 16391, 22997, 23838, 
    25991, 28427, 29640, 30820, 31837, 30318, 28816, 29130, 25310, 21653, 
    18706, 14303, 11524, 6795, 1547, -2104, -5797, -10679, -13493, -17203, 
    -21102, -25005, -26065, -29328, -30430, -31791, -29797, -31079, -29333, 
    -25917, -26697, -21706, -18369, -16663, -10085, -7405, -4258, 432, 4362, 
    10501, 14963, 17649, 19826, 24310, 26013, 28062, 29413, 29772, 30483, 
    30179, 29351, 27371, 25417, 21865, 19379, 14598, 11758, 8383, 3619, 73, 
    -6474, -10419, -13817, -18683, -20399, -24978, -26576, -27885, -28923, 
    -30747, -32128, -30865, -30360, -27578, -24326, -21104, -19684, -14940, 
    -12797, -7348, -2817, -249, 6731, 8402, 12822, 18441, 20247, 23989, 
    25999, 28952, 31145, 31873, 29480, 29568, 29241, 28701, 26129, 23448, 
    20779, 17783, 12567, 7755, 4589, 412, -3616, -9502, -12392, -18638, 
    -21046, -24937, -25962, -28544, -29484, -30709, -30532, -29774, -30139, 
    -28983, -26748, -22207, -20798, -16966, -13230, -8410, -3816, -599, 4707, 
    9407, 14088, 17375, 22208, 22962, 26090, 29961, 30234, 30648, 31058, 
    31560, 29766, 28162, 26853, 22600, 19587, 17338, 13906, 8884, 4025, -95, 
    -4557, -8252, -12398, -16511, -19720, -23603, -25584, -28918, -28868, 
    -30174, -31144, -30565, -29931, -27362, -25738, -21913, -19748, -17158, 
    -13864, -9565, -5506, 67, 5227, 8905, 13436, 16634, 19907, 21497, 25021, 
    28051, 29219, 30584, 32148, 31372, 30359, 28473, 27035, 22575, 20586, 
    18417, 14763, 10022, 5446, -841, -5447, -8485, -11866, -16881, -21376, 
    -23260, -26764, -29223, -28733, -31824, -30134, -30714, -31044, -27169, 
    -26673, -23872, -19977, -16829, -12091, -9633, -3793, 1246, 3539, 6905, 
    11286, 14653, 19405, 22649, 26290, 28917, 30594, 28865, 31009, 29411, 
    29662, 28066, 27432, 23917, 20692, 16646, 13005, 9983, 4741, 1040, -2613, 
    -8669, -12824, -14676, -19005, -22507, -25857, -26726, -30437, -28964, 
    -29633, -29991, -29169, -29943, -25130, -22262, -20296, -17407, -13245, 
    -9995, -5028, -1236, 1737, 7771, 11192, 15771, 18778, 22749, 24363, 
    28008, 31042, 31606, 31437, 30274, 29952, 30038, 25098, 23935, 19731, 
    17283, 12497, 10029, 5303, 1141, -4376, -7397, -11515, -15886, -18583, 
    -23109, -25339, -28180, -28426, -31312, -30877, -30742, -28646, -28514, 
    -26731, -24905, -20885, -18070, -13055, -10033, -6250, -680, 3517, 5825, 
    10939, 14175, 18884, 22777, 23472, 27956, 30742, 30729, 29005, 29582, 
    29469, 27286, 27296, 23447, 22937, 16951, 14183, 11405, 5476, 1090, 
    -2558, -7298, -10462, -15970, -19799, -21780, -25975, -27769, -29339, 
    -31052, -29753, -30895, -29982, -28907, -26665, -24414, -20067, -17731, 
    -15526, -10806, -5093, -466, 2554, 7424, 10632, 16182, 20049, 21755, 
    24806, 26394, 28582, 28930, 31774, 31410, 29760, 27964, 26082, 23345, 
    21599, 19859, 14464, 10426, 6884, 1965, -2769, -7807, -9647, -15705, 
    -18665, -21889, -23328, -28280, -28854, -31524, -32269, -31049, -29546, 
    -28049, -26612, -24218, -21255, -19448, -16358, -9521, -6241, -2424, 
    1558, 5873, 10587, 13486, 18236, 21320, 24897, 26597, 28567, 29201, 
    31952, 30291, 28966, 27994, 26786, 24543, 21798, 18576, 14749, 10588, 
    6744, 1071, -2706, -6176, -11777, -14174, -18347, -22335, -24202, -27798, 
    -27887, -29791, -29699, -30389, -29451, -30807, -28842, -24290, -20998, 
    -19793, -15978, -11958, -7033, -1554, 3599, 4477, 10677, 14205, 18258, 
    22027, 25157, 26266, 30159, 29679, 31480, 31555, 30152, 27773, 27459, 
    23565, 22133, 19003, 14979, 10852, 7165, 3816, -2048, -4818, -10555, 
    -15873, -17217, -20501, -22772, -26297, -27911, -30773, -30581, -30864, 
    -30428, -28670, -26896, -24827, -22736, -18116, -15586, -10411, -6867, 
    -2567, 985, 6040, 11137, 13193, 17317, 21130, 25402, 27187, 27882, 31610, 
    30196, 30396, 31665, 28980, 28887, 25119, 22063, 18221, 16355, 10946, 
    8420, 2032, -1162, -5505, -8572, -13002, -18704, -21540, -23815, -26913, 
    -26733, -28828, -30985, -32123, -31018, -29417, -27877, -24596, -23854, 
    -20491, -15616, -10709, -9300, -3916, 637, 5773, 8997, 14346, 17249, 
    21514, 22717, 26939, 27905, 29348, 29079, 31269, 30613, 28937, 28611, 
    25069, 23917, 18779, 15852, 12296, 7575, 4298, -284, -6025, -10437, 
    -12987, -18372, -20920, -23694, -26021, -28393, -28690, -30014, -30844, 
    -29213, -28998, -26614, -25596, -22648, -18856, -16638, -13052, -9095, 
    -3669, 335, 5100, 9568, 13560, 16802, 20716, 23427, 25648, 27236, 29019, 
    31046, 31803, 31685, 30033, 28032, 25907, 22775, 19169, 17694, 12636, 
    8275, 3586, -1167, -5089, -8599, -13966, -16700, -20507, -24850, -25189, 
    -28261, -29967, -30182, -30243, -30382, -28575, -28906, -26549, -23845, 
    -21197, -16837, -12803, -8921, -3912, -512, 3594, 8316, 12266, 17068, 
    18910, 23501, 24471, 29338, 29764, 29617, 29559, 30222, 29246, 29358, 
    26534, 23057, 19379, 17158, 11776, 8664, 4667, 534, -3821, -8560, -13832, 
    -16829, -19869, -23593, -26120, -27785, -29621, -30561, -32599, -30435, 
    -28734, -28611, -24641, -23210, -19995, -17792, -13398, -9303, -4020, 
    -305, 4039, 7194, 13049, 14768, 18604, 23448, 25577, 28176, 27824, 30115, 
    30253, 31729, 30476, 28106, 25106, 23544, 22053, 16932, 13039, 10232, 
    4389, 1029, -3868, -7870, -13929, -16950, -19716, -21671, -24140, -28339, 
    -28801, -30092, -32245, -30570, -30025, -27981, -25523, -23756, -21440, 
    -19033, -12545, -8796, -4073, -1004, 3375, 9143, 12761, 16391, 19984, 
    21340, 23809, 28698, 29863, 31539, 32141, 30086, 29193, 28519, 25324, 
    23274, 21514, 17713, 12513, 10574, 4510, 816, -2104, -6782, -11558, 
    -16794, -20007, -20860, -25485, -27501, -28536, -29453, -30433, -31126, 
    -30094, -29325, -26609, -23271, -22628, -17004, -14181, -8525, -6867, 
    -774, 2646, 8204, 10758, 16916, 19658, 22858, 25133, 27962, 28860, 31238, 
    31346, 29973, 29655, 27352, 26652, 25033, 21455, 18038, 15037, 11259, 
    4593, 1145, -1360, -7654, -10473, -14877, -18532, -21919, -24281, -27485, 
    -27817, -29543, -29313, -29794, -29060, -29098, -28037, -25673, -22303, 
    -18111, -13687, -11376, -6781, -2639, 2790, 8304, 12743, 16882, 18621, 
    21685, 25672, 26870, 30065, 29128, 30531, 29939, 30507, 28275, 27692, 
    24731, 21049, 17515, 14724, 11583, 8051, 1894, -2209, -5176, -10474, 
    -15959, -17772, -22071, -24680, -28501, -28032, -30405, -30277, -32003, 
    -29575, -28031, -26655, -25613, -22359, -19191, -14708, -10022, -6327, 
    -2276, 1950, 6556, 10785, 15663, 18080, 22173, 25291, 25875, 29819, 
    29464, 31590, 32201, 29370, 28600, 27089, 23625, 21940, 17644, 15811, 
    9620, 6303, 2863, -1076, -6216, -9162, -13718, -18608, -20767, -24647, 
    -26499, -30084, -28748, -28893, -30669, -31511, -30087, -27959, -24681, 
    -22053, -19614, -15343, -10405, -6016, -1537, 1969, 7200, 11466, 13978, 
    16745, 22660, 23153, 27976, 28865, 30473, 31701, 30567, 30802, 28822, 
    25941, 24514, 21163, 20166, 16091, 10547, 7149, 2635, -467, -5438, 
    -10001, -14721, -18444, -22043, -23520, -26932, -28133, -29510, -29789, 
    -31150, -29108, -28290, -27439, -24784, -22424, -18256, -14268, -11016, 
    -8270, -3024, 820, 5874, 11055, 13959, 17325, 19675, 24495, 27606, 27693, 
    30984, 30569, 28981, 30468, 28082, 27728, 25494, 22995, 19152, 17070, 
    11190, 8249, 2784, -298, -4180, -9473, -14309, -17558, -19859, -24255, 
    -27923, -29062, -28797, -30879, -31968, -29947, -29913, -27388, -25865, 
    -23427, -18799, -17336, -11809, -8251, -3215, 90, 4521, 9057, 12917, 
    17031, 21381, 23570, 26268, 29158, 28807, 29407, 30415, 29910, 28861, 
    28077, 26839, 23121, 19758, 16148, 11257, 7040, 3817, -1317, -4555, 
    -10027, -13760, -18177, -20864, -24472, -27230, -27753, -28366, -31457, 
    -31302, -31696, -29688, -26983, -26075, -23486, -19916, -17468, -11931, 
    -8468, -5512, 326, 4408, 9638, 12164, 16985, 21643, 23038, 26289, 28966, 
    30286, 29447, 31123, 31395, 29523, 27343, 25727, 23402, 19610, 15806, 
    12458, 8216, 4520, -1277, -4019, -8186, -12680, -16262, -21000, -23554, 
    -25827, -29477, -29243, -31004, -30066, -30400, -30131, -28408, -26322, 
    -23433, -21524, -17763, -13779, -8635, -4603, -235, 4508, 8940, 11734, 
    17564, 20274, 23709, 26038, 27053, 30202, 29935, 31894, 30353, 29973, 
    27175, 26042, 24799, 18840, 16756, 13222, 9348, 4713, 649, -4054, -8474, 
    -13549, -15162, -21452, -22443, -24162, -28082, -29704, -30462, -31588, 
    -31213, -29311, -27905, -27514, -23149, -19848, -18203, -12005, -9590, 
    -6324, 358, 3282, 9122, 12420, 17154, 19478, 21595, 26317, 26790, 30079, 
    29547, 31310, 30618, 31019, 28507, 26297, 23664, 19916, 18382, 14608, 
    9352, 5566, 923, -3757, -8612, -11200, -16423, -19838, -23938, -26719, 
    -27412, -29561, -30087, -32070, -30488, -28563, -26757, -26353, -24524, 
    -22399, -16402, -14062, -9949, -5221, -2220, 3836, 8610, 11460, 16209, 
    19781, 21949, 26556, 27918, 30726, 29269, 30212, 30063, 29326, 29096, 
    26511, 23129, 21151, 16758, 14078, 8669, 5540, -170, -3671, -6638, 
    -11930, -14976, -19352, -23740, -23701, -26286, -29128, -29736, -30939, 
    -31349, -29007, -29149, -27171, -23244, -20695, -16663, -14652, -9061, 
    -5365, 82, 3097, 7380, 11367, 16985, 19378, 23663, 24397, 26726, 28181, 
    30876, 31770, 30997, 29417, 28338, 26831, 24550, 19465, 17708, 12354, 
    10942, 5571, 1444, -2299, -8458, -12290, -16195, -18981, -23383, -25716, 
    -27302, -30593, -29648, -30060, -30619, -30489, -28845, -27026, -24386, 
    -21770, -18106, -15300, -10456, -6687, -2724, 1813, 5953, 10779, 14977, 
    18843, 22642, 26455, 25485, 28604, 31070, 29407, 30637, 29882, 29640, 
    25663, 24300, 20417, 18306, 13991, 10556, 5984, 3385, -2825, -6771, 
    -9453, -14553, -17799, -20315, -25057, -28613, -30172, -29757, -31470, 
    -31513, -31034, -29402, -26559, -25457, -21852, -18847, -15305, -10232, 
    -5368, -1537, 2471, 5829, 10348, 15164, 17536, 22433, 23629, 27794, 
    29654, 28721, 29235, 30555, 30514, 28725, 27036, 25638, 22483, 18979, 
    15791, 10837, 6816, 3564, -2846, -5159, -10134, -15541, -19744, -21786, 
    -25512, -25919, -28237, -31435, -31703, -29582, -28704, -29881, -25799, 
    -25182, -21358, -18718, -16767, -11190, -6411, -3448, 862, 5556, 10405, 
    14698, 19287, 21061, 24203, 27593, 28574, 29670, 29228, 31996, 29217, 
    28638, 28049, 26749, 22240, 19563, 16112, 10625, 7643, 2584, -2059, 
    -5753, -8892, -15298, -17517, -22311, -24074, -26597, -30215, -30009, 
    -30240, -30251, -31736, -28537, -28199, -26958, -20930, -18580, -14536, 
    -10241, -7522, -3340, 476, 6031, 10053, 14289, 18123, 20712, 24288, 
    26859, 29807, 29695, 30967, 30745, 30108, 29022, 27194, 25802, 22946, 
    18790, 15912, 11771, 6929, 3675, -736, -5125, -9660, -13785, -17764, 
    -20473, -24219, -27409, -28522, -31088, -30616, -29916, -30262, -30880, 
    -25754, -25286, -23781, -20132, -15832, -11582, -6818, -4607, 1186, 3649, 
    9679, 13539, 16580, 19420, 24423, 25591, 28784, 29992, 29507, 30922, 
    31678, 28491, 28340, 25529, 23196, 21026, 15425, 12526, 6723, 4402, -617, 
    -4325, -10874, -12880, -18171, -20664, -24415, -27652, -29711, -30440, 
    -30417, -30571, -30766, -29077, -27352, -25745, -22992, -18416, -15626, 
    -11181, -7111, -3405, -945, 6293, 9076, 13576, 16289, 19761, 24301, 
    26876, 26340, 30835, 29975, 29151, 30034, 28485, 28638, 25634, 22575, 
    19228, 16180, 14066, 9088, 3409, -462, -3802, -8535, -13026, -16131, 
    -19779, -22663, -25333, -27664, -31280, -31139, -29640, -30710, -28468, 
    -27349, -24626, -24277, -20089, -15256, -12865, -9039, -4464, 1251, 4134, 
    8993, 13346, 17814, 19591, 22844, 25907, 27096, 30540, 30644, 31271, 
    29420, 30777, 29310, 26408, 24915, 22115, 16708, 12896, 8148, 4763, 142, 
    -4673, -7562, -12303, -15951, -19644, -23459, -25457, -27812, -29029, 
    -29137, -29755, -30622, -29883, -27110, -25987, -22571, -19421, -16307, 
    -13785, -8557, -4406, -368, 4091, 8277, 13239, 16124, 19762, 21679, 
    25725, 27609, 29806, 28829, 29700, 30873, 30646, 28416, 27941, 23530, 
    20579, 17470, 14184, 10841, 4295, 374, -4636, -8350, -11815, -17119, 
    -18562, -21944, -25503, -29089, -29556, -30365, -31493, -29155, -29929, 
    -27908, -26146, -23833, -21412, -16859, -13695, -8527, -4644, -1731, 
    3531, 6395, 10398, 14981, 19708, 22309, 25276, 27408, 29722, 30209, 
    30841, 30112, 28960, 28714, 26924, 22924, 21672, 17538, 13486, 10480, 
    6558, 1152, -4092, -7428, -11864, -16665, -18885, -23484, -24706, -27725, 
    -29081, -30617, -30528, -30308, -31487, -28156, -27824, -24557, -20703, 
    -17994, -15000, -9403, -5357, -306, 2393, 7385, 11085, 15620, 20313, 
    22773, 26406, 25890, 27340, 30424, 31478, 30496, 30194, 29483, 26560, 
    25021, 21815, 16610, 12983, 10431, 4375, -114, -3029, -6369, -12452, 
    -13933, -17591, -21019, -26045, -27394, -29510, -29308, -30776, -31671, 
    -29414, -28931, -25604, -24813, -21793, -19097, -15505, -10134, -5787, 
    -1603, 3120, 7792, 11436, 14615, 18528, 21624, 24830, 28483, 30218, 
    29254, 31590, 32153, 30246, 29494, 26569, 24615, 22324, 18489, 13895, 
    10306, 6494, 2198, -2288, -7574, -10445, -15850, -18722, -21460, -25104, 
    -26489, -29017, -30122, -30853, -30689, -29788, -28305, -26877, -24287, 
    -22799, -19471, -15271, -11482, -6942, -2810, 2365, 7429, 10774, 14909, 
    18973, 21390, 25873, 27030, 29646, 30691, 31166, 32322, 29005, 29538, 
    26285, 23791, 21082, 18529, 14257, 11167, 6440, 2088, -1412, -6685, 
    -10767, -13540, -19083, -22044, -24704, -25351, -28641, -28541, -30421, 
    -31368, -30761, -27826, -28568, -24635, -21092, -18521, -16174, -10120, 
    -7047, -4143, 1644, 6055, 10840, 14945, 17873, 19918, 24750, 28310, 
    29753, 28920, 32335, 30990, 30813, 28598, 27296, 24464, 23199, 17793, 
    13977, 10487, 7255, 2418, -886, -4889, -10916, -13813, -17775, -20227, 
    -22800, -28114, -29665, -29028, -31221, -30123, -29164, -29780, -27370, 
    -24546, -21364, -18337, -14170, -12646, -7152, -3171, 1921, 5390, 10640, 
    14815, 17573, 20647, 25228, 27608, 27541, 30751, 31302, 30261, 28856, 
    29280, 27804, 26265, 23953, 19252, 15509, 12187, 8812, 1858, -968, -4213, 
    -9256, -12863, -18419, -20163, -24183, -25650, -27582, -31584, -30788, 
    -31237, -31476, -29082, -26614, -25010, -22791, -19012, -15384, -13164, 
    -7560, -3261, 1645, 6771, 10542, 12217, 17278, 21021, 22814, 24602, 
    29356, 28967, 31190, 31258, 31847, 29134, 26221, 25900, 22356, 19591, 
    16288, 10928, 6323, 4690, -1003, -3342, -9931, -13199, -16333, -20232, 
    -23524, -25589, -27945, -30454, -30281, -31736, -30320, -30953, -28034, 
    -25359, -22240, -20253, -15743, -12138, -6631, -4981, 87, 6352, 10021, 
    13454, 16877, 21803, 22444, 27078, 28013, 29619, 31043, 30569, 31912, 
    30947, 28177, 25709, 22551, 19985, 16206, 12832, 7776, 4842, 775, -5551, 
    -10754, -11902, -17279, -20515, -23880, -26522, -27680, -28876, -29176, 
    -30048, -30009, -30183, -27942, -25618, -23788, -19623, -16077, -12447, 
    -9840, -3843, 220, 3458, 8855, 12855, 16423, 20342, 24594, 24998, 28010, 
    28275, 31877, 29789, 30298, 29193, 29710, 26236, 23096, 20821, 16845, 
    12963, 8134, 4433, 1120, -3797, -9096, -12693, -15886, -19049, -24597, 
    -25671, -28036, -30993, -30178, -31283, -31762, -29758, -29405, -27400, 
    -23465, -20953, -18301, -12017, -8183, -4089, -563, 4544, 7785, 12546, 
    15115, 18916, 22555, 24368, 27505, 28579, 30540, 30973, 29550, 29084, 
    27171, 26040, 23222, 19837, 16323, 13137, 9714, 4619, 731, -3256, -8233, 
    -11295, -15376, -18325, -23292, -25147, -28545, -30337, -31001, -31600, 
    -29158, -28889, -29672, -25571, -23633, -19941, -16194, -14428, -9572, 
    -5712, -779, 3336, 8725, 12546, 15618, 18966, 24509, 26158, 27027, 29199, 
    30614, 31628, 31039, 30104, 28608, 26886, 22793, 21424, 17273, 13991, 
    10942, 5662, 1020, -3495, -6717, -10407, -14732, -20597, -22226, -25067, 
    -27303, -28004, -30244, -30276, -29295, -30953, -27498, -27612, -24519, 
    -21315, -17826, -12810, -8513, -5622, -1207, 3277, 8648, 12073, 16252, 
    18753, 22609, 24203, 27957, 27789, 31425, 30849, 30056, 28526, 27721, 
    26765, 25662, 22128, 18776, 14315, 10223, 6521, 2399, -2546, -5697, 
    -11852, -15797, -19782, -21533, -24934, -27587, -27939, -29872, -30611, 
    -29763, -30535, -29024, -26816, -24036, -21525, -17894, -15033, -10684, 
    -7025, -2028, 2523, 6572, 12285, 14344, 18294, 23805, 25923, 28602, 
    28355, 30195, 31098, 31798, 29151, 29814, 28002, 25043, 22876, 17525, 
    15754, 11210, 5906, 2019, -3368, -7030, -11169, -15288, -19126, -22679, 
    -25507, -27450, -28852, -30395, -31588, -29144, -30117, -28875, -26505, 
    -25824, -21037, -19146, -14957, -11357, -7938, -2380, 3749, 6188, 10766, 
    14924, 17968, 21854, 23979, 27554, 28699, 29521, 31726, 31895, 31279, 
    28667, 27352, 25335, 23214, 18240, 15348, 12093, 8669, 2733, -1399, 
    -6032, -10157, -14813, -18242, -22668, -25321, -27294, -30215, -28489, 
    -31680, -32150, -30045, -28663, -27813, -26441, -23547, -17370, -14720, 
    -11244, -5730, -2353, 2077, 6356, 11086, 15628, 18608, 21319, 23799, 
    26557, 28754, 28827, 29773, 31418, 31718, 29565, 27030, 24589, 22850, 
    18300, 15090, 11855, 6433, 2113, -1714, -6107, -10495, -13867, -18149, 
    -22358, -23535, -26277, -29029, -28699, -29270, -29992, -30635, -28778, 
    -27657, -26324, -22042, -19895, -16388, -11431, -7975, -3510, 1662, 4683, 
    10474, 14413, 17185, 20292, 23972, 27064, 26773, 28937, 30003, 30038, 
    31167, 29103, 27719, 25627, 22696, 19134, 15431, 12179, 6352, 4305, 232, 
    -4695, -9764, -13038, -17052, -21635, -23240, -25030, -28729, -30374, 
    -31304, -31764, -30884, -30376, -26935, -25717, -22301, -19899, -16055, 
    -12704, -8810, -2138, 2661, 6481, 10354, 14868, 17592, 19802, 23379, 
    26292, 28636, 30324, 31131, 30344, 30401, 29460, 26966, 25316, 21540, 
    19596, 16094, 13024, 6882, 4194, -1477, -4983, -9648, -11862, -16360, 
    -18982, -23629, -26905, -27223, -28672, -29433, -30242, -29611, -30077, 
    -29462, -26888, -24105, -19755, -15918, -11453, -8542, -4359, -644, 6008, 
    8879, 11587, 17590, 21112, 23931, 26424, 29462, 30887, 31012, 31983, 
    29873, 28884, 28716, 24718, 23901, 20553, 16389, 13559, 8067, 4118, 
    -1045, -4773, -9040, -13007, -15479, -21239, -24279, -26146, -26748, 
    -29675, -31002, -32286, -29023, -30708, -27821, -25203, -24325, -19924, 
    -15443, -13572, -8464, -4785, 1132, 4157, 8544, 13925, 16661, 20566, 
    23122, 25805, 27778, 29050, 31321, 31112, 30749, 29179, 29066, 25170, 
    24072, 21185, 16989, 14532, 9659, 4844, -68, -3331, -9321, -13320, 
    -16865, -18869, -22165, -25634, -28721, -29064, -30333, -29498, -29048, 
    -29186, -28534, -25926, -24368, -19959, -18595, -13865, -8112, -4552, 
    476, 4291, 7755, 12928, 17546, 21448, 23569, 25227, 27534, 28344, 30101, 
    31049, 29650, 29099, 28724, 25794, 22710, 20644, 17337, 14350, 8783, 
    5755, 78, -4833, -8450, -10919, -15972, -20015, -22765, -24080, -27087, 
    -28177, -30988, -31546, -29944, -30186, -29167, -26523, -22585, -21953, 
    -16253, -14772, -8830, -6501, -1196, 3668, 7470, 11884, 17562, 18146, 
    22659, 25925, 26042, 27889, 31316, 31053, 32327, 28914, 29447, 26382, 
    23512, 21167, 16445, 14378, 8742, 6511, 1443, -2862, -7207, -12783, 
    -15032, -18964, -24424, -25049, -27434, -29216, -29657, -31957, -31478, 
    -31117, -28931, -26686, -22680, -20869, -17725, -14537, -10053, -6965, 
    -1226, 1935, 7623, 11706, 15008, 18696, 23047, 25162, 28613, 29864, 
    30592, 30164, 29926, 30613, 28035, 27816, 23581, 20978, 17109, 14030, 
    9874, 6270, 2568, -4268, -6197, -9753, -13982, -19511, -22665, -25109, 
    -27739, -28967, -29698, -30753, -30671, -30902, -28127, -27145, -23208, 
    -22570, -18609, -13310, -9956, -5538, -1962, 1292, 6967, 11378, 15068, 
    18271, 23285, 24938, 27749, 29028, 29621, 30557, 29190, 29845, 29292, 
    26216, 24673, 20331, 17957, 15094, 9616, 6317, 2662, -2964, -5291, 
    -10364, -15499, -19951, -20787, -25773, -26779, -28565, -29867, -30369, 
    -31687, -29559, -28068, -27054, -25007, -21493, -17706, -13927, -10486, 
    -5592, -1934, 2340, 6296, 9838, 13849, 18789, 21518, 24651, 26542, 27007, 
    30665, 30703, 31655, 28734, 29329, 25994, 24516, 23149, 18634, 13918, 
    11824, 6377, 3401, -2819, -5494, -10999, -14958, -17972, -21543, -24563, 
    -27226, -28191, -29125, -30116, -30933, -30177, -29545, -27674, -25554, 
    -21614, -18909, -15402, -11205, -7533, -3081, 1354, 5373, 11295, 14979, 
    16983, 22617, 22989, 26607, 28598, 30535, 31625, 29816, 28806, 29499, 
    29133, 25163, 20709, 18660, 16428, 12260, 6265, 2430, -202, -5471, -9309, 
    -14201, -18000, -21227, -24036, -27543, -30046, -29938, -30831, -31799, 
    -29729, -29837, -26830, -25440, -22871, -17990, -14658, -11399, -8360, 
    -2867, 677, 5187, 10598, 12677, 17222, 21490, 23238, 25228, 29825, 29681, 
    29088, 30058, 29233, 30388, 27837, 25282, 21482, 19697, 15726, 12770, 
    9001, 3891, -74, -4377, -10308, -12479, -17629, -21741, -23820, -26050, 
    -28172, -30451, -30314, -30739, -29811, -29923, -27472, -25622, -21701, 
    -21002, -14608, -12691, -7535, -2503, 1156, 3904, 9216, 13209, 16655, 
    20897, 22543, 25650, 26883, 29088, 30559, 30368, 30432, 29228, 27828, 
    25586, 24113, 19543, 15856, 11634, 7892, 3196, 496, -3247, -9685, -13418, 
    -17880, -21785, -22846, -27391, -27951, -30706, -28964, -31047, -30372, 
    -28571, -27252, -25163, -23719, -20380, -17144, -12387, -7520, -3933, 
    1846, 5923, 7440, 13103, 17054, 21555, 24010, 27435, 26530, 28663, 30867, 
    30634, 29404, 30415, 28358, 25981, 22965, 19261, 16207, 12879, 8103, 
    4342, -831, -4921, -8644, -13042, -16439, -22114, -23995, -26203, -29134, 
    -29672, -30057, -29894, -29756, -28594, -28070, -25278, -21901, -20143, 
    -16619, -12882, -8954, -3444, -758, 3252, 9663, 13785, 16769, 19553, 
    23059, 24101, 26863, 29012, 32076, 30749, 32083, 30278, 28989, 24201, 
    22899, 20095, 16817, 13716, 8877, 3720, -67, -2785, -9834, -11590, 
    -16933, -19638, -21780, -26212, -28812, -28555, -30815, -29198, -31066, 
    -29944, -26621, -26118, -21883, -20755, -17159, -14057, -10227, -5206, 
    -395, 4983, 7819, 12445, 15776, 20752, 22430, 25564, 28674, 30779, 29832, 
    30229, 30205, 30521, 30012, 25583, 24398, 21842, 17355, 12882, 8597, 
    4530, 946, -3049, -7915, -12244, -15373, -19488, -23505, -26809, -26796, 
    -30721, -29490, -31403, -31519, -29177, -28790, -25942, -25020, -20016, 
    -17380, -13921, -9460, -6117, -2190, 2128, 9039, 11816, 14409, 19732, 
    21463, 25641, 26923, 29631, 30338, 31180, 30177, 29790, 28523, 27128, 
    25722, 20746, 17554, 14601, 9348, 7357, 1251, -2814, -7831, -10591, 
    -16234, -18432, -22349, -25635, -27607, -28521, -29049, -31887, -29785, 
    -29087, -29527, -26647, -23559, -22212, -18956, -15594, -8923, -6432, 
    -1590, 1970, 6450, 11993, 15517, 19050, 22355, 25464, 26946, 30176, 
    29882, 29162, 30923, 30317, 27614, 26301, 24550, 20497, 19125, 14571, 
    9349, 6142, 1248, -3589, -6619, -9857, -15985, -19842, -21472, -25564, 
    -27410, -29427, -31647, -31260, -29909, -31328, -30144, -26155, -23525, 
    -20568, -18155, -13372, -10229, -5306, -668, 1637, 7789, 11486, 14446, 
    16944, 22355, 25286, 27176, 28296, 30836, 30748, 30386, 30457, 27575, 
    27447, 24989, 21389, 19374, 14609, 10427, 6958, 2629, -3932, -6832, 
    -11361, -14298, -18091, -21659, -24652, -26689, -30223, -29667, -30690, 
    -30190, -29560, -28883, -26831, -25332, -22900, -17296, -14279, -11939, 
    -6546, -1621, 2038, 7187, 11663, 13815, 19782, 20992, 25537, 28568, 
    29944, 29952, 29789, 31586, 30351, 30222, 26297, 24646, 20633, 19919, 
    15445, 11429, 5484, 2025, -2294, -5162, -11271, -16046, -18380, -23073, 
    -24093, -25920, -28579, -30315, -31569, -31974, -30243, -29464, -28868, 
    -24309, -21428, -19220, -15398, -9620, -7371, -2684, 1866, 6979, 10995, 
    14487, 17124, 21011, 23486, 27995, 28620, 29483, 31789, 30631, 29340, 
    29137, 27070, 24543, 21896, 19347, 16805, 10830, 6768, 3599, -2276, 
    -4870, -9535, -14340, -18212, -21654, -24971, -27550, -29303, -30145, 
    -31805, -31431, -29254, -28748, -26057, -25336, -23308, -18331, -16665, 
    -11912, -7067, -2297, 826, 6006, 10483, 13815, 18473, 21032, 23051, 
    26704, 27068, 30342, 31145, 31524, 30646, 28569, 27952, 24955, 23006, 
    19008, 15035, 12777, 7562, 1978, -906, -7334, -9534, -12931, -18481, 
    -19612, -23574, -26834, -27730, -28967, -30347, -31264, -29778, -30132, 
    -27353, -24894, -23349, -19367, -16670, -12404, -6445, -3777, 2386, 4907, 
    8866, 15078, 17652, 21347, 24658, 26622, 27391, 28651, 30650, 31277, 
    30032, 28815, 29451, 24610, 22575, 20526, 17783, 11238, 7338, 3604, -700, 
    -4079, -8561, -12152, -17576, -20854, -22742, -26431, -28612, -30609, 
    -30285, -31530, -31554, -30244, -26421, -24726, -21907, -19690, -14762, 
    -12509, -7740, -2969, 494, 5104, 10967, 13101, 16920, 21430, 22407, 
    26195, 28455, 29308, 31375, 31786, 29243, 28599, 28623, 25284, 24206, 
    18967, 17322, 12567, 7147, 2866, -846, -4270, -8168, -12867, -17612, 
    -19132, -24251, -26263, -28533, -28631, -30746, -30649, -30305, -29434, 
    -28044, -26538, -21904, -19308, -17536, -13736, -9211, -3593, 786, 5356, 
    8321, 12420, 15634, 18928, 22129, 25424, 28641, 29890, 31769, 31753, 
    31465, 30860, 28404, 26158, 24670, 20757, 15918, 12844, 9925, 4412, -527, 
    -2449, -9495, -13097, -15613, -19701, -21691, -25498, -27995, -29461, 
    -30946, -30802, -29325, -29134, -28362, -25240, -24369, -19703, -16655, 
    -12397, -7974, -3939, -1443, 3664, 9877, 11950, 17860, 19819, 23958, 
    26563, 28097, 31319, 30165, 29807, 30464, 28623, 28916, 25473, 22968, 
    20327, 17628, 13640, 8687, 4158, -778, -3117, -9040, -10999, -16555, 
    -18725, -22999, -26972, -28425, -29340, -30856, -30192, -30172, -29732, 
    -28657, -25989, -24484, -21195, -17662, -14216, -9150, -5402, -1011, 
    4491, 8047, 12450, 16157, 20875, 21939, 24597, 28584, 28571, 30688, 
    31015, 30347, 31172, 28040, 25579, 23074, 20950, 17690, 13944, 9177, 
    4782, 907, -3040, -8569, -10247, -15797, -20074, -22907, -26539, -27710, 
    -30668, -30379, -31362, -29677, -28919, -30164, -26764, -23648, -20810, 
    -16858, -14470, -10254, -5977, -1941, 4169, 6491, 11875, 15727, 20785, 
    22551, 26383, 28934, 30066, 31176, 31538, 29846, 29526, 29272, 27800, 
    24545, 20122, 18644, 13277, 11250, 5476, 1938, -3215, -7975, -12297, 
    -16985, -19584, -22569, -24296, -25975, -27698, -30991, -32481, -31041, 
    -30217, -29384, -26649, -24549, -20348, -17476, -13566, -9372, -5890, 
    -2101, 2980, 6577, 9949, 15277, 17205, 23899, 26555, 27784, 29932, 30073, 
    29991, 29426, 29428, 29631, 26800, 24297, 21669, 16785, 14319, 11126, 
    6766, 996, -3796, -6432, -11103, -15448, -18961, -22417, -24628, -27919, 
    -29673, -32014, -30803, -30160, -30656, -27480, -26864, -24763, -21306, 
    -17221, -13700, -9941, -7883, -3561, 1232, 5033, 10288, 14638, 18852, 
    21619, 25705, 27799, 28364, 30858, 30568, 30171, 29424, 28513, 27772, 
    25661, 22088, 19262, 15334, 10948, 7063, 2006, -1471, -5944, -11614, 
    -15144, -18756, -21374, -25080, -28177, -28064, -29321, -30479, -29636, 
    -30287, -28506, -26433, -24464, -22270, -19626, -14037, -10478, -8276, 
    -2087, 672, 4711, 10415, 14111, 18249, 22071, 24741, 27723, 28178, 28543, 
    30114, 30192, 31527, 30163, 28194, 23645, 21682, 17903, 15712, 12291, 
    8442, 2070, -2874, -5706, -11851, -14961, -17710, -22356, -25151, -26285, 
    -28453, -30087, -31437, -29951, -30522, -30337, -28059, -24879, -22604, 
    -18651, -16099, -10326, -7945, -2353, 1515, 5430, 8747, 13326, 18405, 
    22007, 24605, 25616, 28935, 28669, 29986, 30305, 29976, 28224, 28207, 
    26634, 21602, 20885, 15192, 11142, 8342, 2226, -1552, -4679, -10715, 
    -13024, -18363, -20782, -23892, -26630, -28458, -29146, -30379, -30854, 
    -29083, -29693, -26998, -25300, -22728, -18788, -16040, -10071, -8231, 
    -4508, 957, 4060, 11110, 13503, 16254, 20803, 25500, 25484, 28350, 30880, 
    29928, 31428, 30643, 28644, 28887, 25124, 22334, 19757, 16493, 13766, 
    8267, 4123, -113, -6630, -10476, -13423, -17643, -20771, -23868, -25234, 
    -29208, -28594, -32028, -31286, -30980, -29601, -27618, -24470, -22954, 
    -20637, -14895, -12431, -9293, -2900, 890, 5758, 9562, 11460, 16691, 
    20517, 23671, 25943, 27111, 29485, 29251, 31499, 31045, 29343, 28053, 
    26050, 23662, 20138, 15785, 13216, 8394, 4271, 171, -6199, -8057, -13989, 
    -15404, -20738, -23888, -24269, -29790, -28713, -29715, -29791, -30823, 
    -29844, -27425, -26335, -24749, -18658, -15706, -11985, -8933, -4680, 
    -398, 3648, 9314, 12554, 16976, 21614, 23291, 25877, 27369, 29069, 31397, 
    29691, 31016, 30487, 27288, 26387, 22193, 21381, 16020, 12000, 9463, 
    5286, 1507, -4620, -8216, -12040, -15688, -20843, -23929, -25658, -28038, 
    -29131, -31194, -31230, -30591, -29546, -28747, -26850, -24703, -20763, 
    -17264, -12580, -9689, -4244, -1466, 4652, 8513, 12068, 15948, 20105, 
    22539, 25738, 26869, 30492, 30527, 32059, 29235, 28754, 28717, 27070, 
    23933, 21023, 16424, 13168, 8379, 5278, 1527, -2594, -8026, -12575, 
    -14870, -19282, -22741, -25166, -27606, -28487, -30499, -30692, -30709, 
    -30270, -29569, -26530, -24538, -21765, -16073, -14137, -10861, -6702, 
    -1173, 4285, 8650, 11058, 14905, 17844, 22561, 26393, 28133, 28052, 
    30679, 31462, 30966, 30500, 29374, 26998, 25313, 20688, 17079, 14811, 
    8833, 4255, 2208, -3383, -7139, -11679, -15546, -18755, -23723, -24476, 
    -28069, -28486, -30820, -30890, -31291, -29861, -28427, -26014, -24105, 
    -21999, -18573, -13566, -10753, -5217, -2598, 3754, 6979, 12312, 14201, 
    18707, 22320, 25569, 27721, 29460, 29436, 29753, 30039, 29507, 28706, 
    28205, 24784, 21791, 17173, 13763, 10097, 6120, 859, -2758, -6849, 
    -11496, -15657, -19840, -21863, -26253, -27144, -28728, -30951, -28975, 
    -31946, -30380, -27854, -27916, -24591, -21192, -18814, -15829, -9376, 
    -5474, -1921, 3219, 5960, 11923, 15110, 18468, 22676, 23508, 28341, 
    28729, 30273, 32251, 31140, 28914, 29718, 26962, 24241, 22705, 18593, 
    14682, 10859, 4676, 1970, -2787, -5771, -10456, -15560, -18735, -22227, 
    -23867, -27300, -27845, -31660, -31040, -30131, -31004, -28599, -27534, 
    -24435, -20549, -19398, -14463, -11661, -5909, -3038, 2357, 6622, 9803, 
    13491, 17505, 22215, 26208, 27133, 29081, 29153, 30096, 30834, 29630, 
    29959, 27681, 26058, 21261, 19331, 13350, 10631, 6044, 1379, -2753, 
    -5710, -11435, -13968, -19071, -22041, -24632, -27304, -29008, -30855, 
    -30174, -31636, -31080, -30160, -27341, -23498, -21481, -17930, -13350, 
    -11712, -5659, -3526, 2392, 7338, 10011, 14304, 17479, 22298, 22897, 
    26805, 28439, 29783, 30687, 31111, 29932, 29478, 27219, 25753, 22597, 
    19989, 14500, 10687, 7845, 2987, -2246, -6373, -9075, -15990, -17037, 
    -22398, -24958, -27841, -28440, -30934, -31653, -32410, -31773, -27908, 
    -26702, -23845, -20908, -19193, -15960, -12531, -7165, -2450, 1783, 5948, 
    8918, 12615, 17518, 21921, 25229, 26842, 27771, 31179, 31276, 31089, 
    30394, 28602, 27816, 25553, 21258, 20095, 16079, 12549, 7055, 1955, -850, 
    -4432, -10566, -14484, -16102, -21003, -24847, -25991, -29664, -29109, 
    -30024, -30021, -30390, -28194, -27637, -25167, -22600, -18695, -17006, 
    -11242, -7582, -4790, -777, 5303, 8158, 14932, 17700, 21806, 24361, 
    25886, 29219, 30295, 29008, 29873, 30559, 29103, 26246, 26082, 23623, 
    19749, 16390, 12116, 7363, 2383, -243, -4750, -10342, -12695, -16998, 
    -20979, -23449, -25700, -29108, -29599, -31393, -31729, -30757, -30914, 
    -27459, -24593, -23733, -19698, -15986, -12008, -8183, -4969, 32, 4714, 
    7671, 13420, 16208, 20202, 23329, 25580, 27915, 29993, 30469, 30897, 
    30963, 29047, 27735, 27287, 23196, 18866, 16824, 12737, 8571, 3423, 979, 
    -4881, -9893, -12389, -17873, -20699, -22859, -27403, -27429, -31038, 
    -29521, -31928, -30750, -30034, -27432, -24741, -23333, -21623, -15636, 
    -12238, -8691, -5831, -1260, 4534, 7948, 12062, 15721, 19909, 24265, 
    24200, 26630, 30975, 31599, 32150, 30788, 28827, 28308, 25001, 24018, 
    19779, 16359, 12530, 9073, 4336, 326, -3368, -8967, -12207, -16893, 
    -19667, -22720, -25858, -27753, -29930, -31035, -30906, -29746, -30146, 
    -26386, -24785, -23394, -20564, -17008, -12592, -9886, -5110, 53, 4400, 
    7935, 13530, 17673, 19233, 22868, 25371, 28572, 29075, 30155, 31475, 
    30837, 30868, 27738, 26432, 24692, 19686, 17221, 12595, 9850, 5179, 1464, 
    -4654, -8877, -12318, -15324, -19053, -23044, -24059, -26603, -28457, 
    -28607, -30755, -30743, -30496, -28419, -25595, -24695, -20039, -18893, 
    -13858, -8902, -5649, 467, 2942, 8255, 11338, 15993, 18009, 23796, 26826, 
    27735, 29549, 29929, 31390, 32162, 29143, 28403, 28267, 23325, 20061, 
    18398, 15037, 10144, 5045, 2370, -3085, -6615, -11802, -15270, -18809, 
    -23651, -24279, -26694, -29193, -31021, -31770, -29346, -28906, -27750, 
    -25660, -24997, -22758, -17759, -12394, -8629, -6721, -1446, 2858, 6193, 
    12652, 15657, 19268, 22519, 24260, 25982, 27818, 28898, 29804, 30316, 
    29287, 27844, 25353, 23926, 22004, 18390, 14643, 10475, 5677, 2462, 
    -2408, -6901, -10382, -15956, -19185, -22164, -25454, -26906, -28339, 
    -29566, -31286, -30455, -30083, -29059, -27200, -25549, -20971, -17876, 
    -15474, -10110, -5526, -3033, 3797, 7670, 11997, 15757, 18741, 23615, 
    24404, 26321, 28633, 30252, 31633, 30474, 31302, 30238, 26710, 24810, 
    23032, 17470, 13425, 11237, 4850, 1459, -2676, -7545, -10674, -14372, 
    -18836, -20232, -24922, -26334, -28889, -30990, -30767, -30452, -31089, 
    -29422, -27226, -24444, -22244, -16654, -14362, -11247, -6948, -1839, 
    2581, 7643, 11131, 15399, 17193, 21653, 24564, 27632, 27803, 29586, 
    30785, 31007, 29269, 30221, 28254, 24028, 21162, 17521, 15224, 10845, 
    6789, 1645, -3226, -6658, -11170, -16137, -17278, -20549, -24543, -26886, 
    -29013, -28774, -29779, -30978, -28671, -27964, -28518, -24069, -21342, 
    -19643, -14249, -9879, -8545, -4295, 676, 6938, 9290, 15253, 18695, 
    20458, 24731, 26698, 28428, 30767, 30507, 29859, 31957, 29220, 25887, 
    26236, 22403, 19431, 15952, 11149, 8739, 1872, -2225, -6457, -9455, 
    -15741, -17864, -20457, -23706, -26640, -28426, -29276, -30165, -29864, 
    -29027, -28210, -25818, -25455, -23098, -19063, -16072, -11247, -7399, 
    -1817, 1476, 7234, 10421, 12751, 18654, 20807, 23644, 27497, 29432, 
    30219, 30236, 32411, 30457, 29953, 28071, 25774, 22484, 18082, 14716, 
    12655, 8467, 4677, -619, -5905, -9777, -14207, -17619, -21595, -24465, 
    -27314, -29393, -29804, -30979, -30043, -30845, -29255, -27508, -25026, 
    -23032, -19499, -14369, -12609, -7445, -3783, 1269, 5545, 8570, 12380, 
    18609, 21226, 24088, 26711, 27221, 29875, 31370, 29677, 31433, 28489, 
    27126, 26178, 23089, 20142, 16693, 13133, 7377, 3483, -705, -5494, -9728, 
    -11969, -17011, -20578, -23578, -24695, -26586, -30200, -29772, -31461, 
    -30209, -29103, -27223, -25470, -23426, -19340, -17021, -11658, -7852, 
    -2956, 1106, 5714, 9692, 12151, 17176, 20250, 24105, 25947, 28510, 30211, 
    30917, 30465, 29605, 31078, 26381, 26147, 24275, 18646, 16072, 13549, 
    7290, 4301, 618, -4742, -8802, -11955, -16584, -21570, -22502, -26808, 
    -28495, -29349, -30134, -31243, -29874, -28467, -28436, -25694, -24623, 
    -21902, -16843, -11562, -7450, -3584, 663, 4156, 8290, 12894, 16089, 
    20151, 23268, 25981, 27691, 28615, 30190, 30831, 30315, 29695, 28003, 
    26450, 22248, 19549, 15448, 13733, 8712, 4178, -1318, -4054, -7705, 
    -11483, -16042, -20162, -22349, -25881, -28807, -28043, -30350, -30177, 
    -31536, -29236, -28706, -26829, -22644, -19778, -16199, -12868, -9627, 
    -5299, -576, 4275, 8259, 11556, 16024, 20449, 22625, 26351, 28398, 28939, 
    31358, 31648, 30769, 29573, 28069, 26575, 24128, 21152, 17521, 13449, 
    8598, 6100, 2398, -3188, -8153, -12167, -17690, -18853, -23200, -25249, 
    -28822, -30335, -29991, -29958, -30541, -31490, -27759, -25092, -22844, 
    -20538, -17064, -11708, -10238, -4972, -700, 3159, 8265, 11454, 15812, 
    20662, 24182, 24458, 27681, 29197, 31581, 30422, 29944, 29589, 28679, 
    26768, 23376, 22188, 18238, 12960, 9292, 6185, 663, -4109, -7346, -12781, 
    -16763, -19673, -21952, -23959, -27265, -29881, -31177, -28998, -30496, 
    -30996, -28238, -26557, -22940, -22338, -17437, -14089, -9295, -6854, 
    -994, 3100, 8011, 12656, 15083, 20619, 22098, 25847, 26888, 28179, 30240, 
    32060, 32204, 29399, 28200, 25661, 25250, 21664, 18907, 13086, 11443, 
    5664, 2172, -2632, -8442, -12338, -15564, -19261, -22340, -25216, -28130, 
    -27829, -30607, -30349, -31174, -30783, -27264, -25432, -23762, -23097, 
    -17937, -15618, -9571, -5974, -2350, 3143, 6262, 11555, 14453, 18365, 
    22571, 24846, 26516, 27727, 29864, 30000, 30954, 30229, 30431, 27171, 
    25140, 22096, 18358, 14811, 10305, 4886, 2811, -1970, -6279, -11730, 
    -14762, -18018, -22100, -23898, -25650, -29828, -29566, -30708, -30501, 
    -29895, -29835, -25616, -24904, -22342, -19188, -14814, -11779, -7009, 
    -2148, 1848, 6127, 9694, 15234, 17264, 22406, 25540, 26413, 28683, 28809, 
    29598, 30729, 31320, 30005, 27436, 25285, 22531, 18265, 14487, 11011, 
    6553, 1164, -3411, -6613, -11933, -14897, -18086, -21996, -25689, -26699, 
    -27986, -30806, -29322, -30921, -30127, -29683, -25806, -24790, -23582, 
    -17725, -15210, -12186, -8668, -3304, 1499, 6271, 10450, 14785, 19044, 
    22089, 23376, 27428, 28284, 28972, 30237, 29872, 31691, 30300, 28511, 
    25738, 22758, 18226, 16071, 10290, 6803, 3812, -1395, -5022, -10793, 
    -14475, -17924, -21755, -23911, -27025, -27988, -30096, -31566, -30694, 
    -29617, -29482, -28399, -25086, -21584, -19891, -16280, -12383, -7979, 
    -4330, 145, 5259, 9383, 13009, 16328, 22838, 23222, 26757, 28749, 31380, 
    30254, 29987, 29500, 27863, 26293, 24568, 21200, 20097, 15636, 10769, 
    7192, 2938, -433, -5177, -9974, -14394, -17094, -20335, -23501, -26852, 
    -28137, -29625, -31601, -31223, -30553, -30440, -27527, -25876, -23202, 
    -21232, -16534, -12041, -8973, -3531, 2628, 5379, 9375, 14506, 17748, 
    19254, 23892, 26389, 27869, 29338, 31394, 31260, 30613, 29359, 27111, 
    25338, 23973, 20166, 16527, 11445, 6756, 3968, -1438, -4552, -8829, 
    -15082, -17650, -20592, -24669, -25564, -28025, -30519, -30539, -29340, 
    -29869, -28231, -26704, -25242, -23966, -21359, -15137, -11860, -8501, 
    -3663, -1, 4340, 10018, 12735, 16182, 20657, 23568, 27486, 28572, 28313, 
    31113, 29272, 29489, 29180, 26915, 26618, 24314, 20295, 14842, 11292, 
    7184, 4154, -183, -5892, -8433, -14091, -16272, -18891, -22565, -26631, 
    -27960, -27781, -29797, -29483, -29849, -30764, -27823, -25120, -24053, 
    -19871, -17903, -13150, -7831, -3465, 935, 5916, 8179, 12554, 16777, 
    19466, 24735, 26193, 28543, 28384, 31878, 30723, 30395, 31259, 26902, 
    26555, 24285, 19117, 15560, 12361, 9736, 3706, 134, -3888, -8375, -11986, 
    -16350, -20443, -23000, -25497, -26960, -29053, -30773, -31122, -31740, 
    -29800, -28403, -26015, -23341, -20525, -16583, -13972, -9166, -3306, 
    -1466, 4855, 7791, 11476, 15890, 19330, 23079, 24540, 28801, 29551, 
    30560, 31788, 31206, 29599, 29211, 25016, 24876, 20253, 17055, 12695, 
    9735, 4771, 1135, -3450, -7867, -10943, -15271, -20161, -23670, -25163, 
    -28987, -29133, -31137, -32195, -31792, -29431, -29056, -26063, -24746, 
    -20349, -17189, -13559, -8765, -5461, 745, 4291, 7778, 11524, 16455, 
    20018, 21171, 25283, 28199, 28775, 30659, 30928, 31973, 29105, 28259, 
    25233, 25363, 20607, 18468, 14309, 10001, 4101, -414, -3475, -7397, 
    -11859, -15520, -20935, -23057, -25077, -28292, -29721, -31309, -31105, 
    -29433, -30337, -29746, -26439, -24415, -22559, -18317, -13348, -9993, 
    -5175, -1838, 3587, 6994, 11172, 13748, 17371, 22223, 26273, 27128, 
    28181, 30712, 29586, 29430, 29037, 26853, 27212, 24104, 21497, 18809, 
    13170, 8540, 4661, 2557, -4421, -6925, -10039, -14884, -19324, -22063, 
    -26032, -28297, -30462, -29768, -31133, -30118, -30057, -28524, -27493, 
    -23810, -20832, -17145, -14571, -11576, -5527, -704, 3122, 6732, 10396, 
    15605, 20280, 21424, 24065, 26880, 29192, 29712, 32377, 30411, 31209, 
    30427, 26461, 24701, 21805, 19458, 13979, 11008, 5390, 1260, -824, -6562, 
    -10783, -14632, -18993, -22228, -23881, -25959, -28265, -30506, -31739, 
    -31154, -29618, -28477, -27354, -24762, -22893, -19785, -14434, -9957, 
    -5575, -2610, 2804, 4960, 11362, 15546, 18542, 22042, 24787, 26551, 
    28112, 30116, 29313, 31781, 30230, 29148, 27801, 24159, 20359, 18420, 
    13359, 9649, 7956, 2702, -3452, -5748, -10484, -14595, -17368, -22499, 
    -25151, -27744, -28771, -29592, -32012, -31352, -30888, -29645, -26831, 
    -25032, -22147, -19119, -16363, -11851, -6461, -3048, 73, 7579, 10846, 
    13983, 18316, 19955, 23462, 27261, 28704, 30610, 30012, 30943, 30473, 
    28116, 27583, 25841, 21722, 17676, 15608, 10341, 7471, 2550, -1686, 
    -6827, -9310, -14531, -18090, -20368, -24244, -25237, -27207, -29430, 
    -30716, -31425, -30560, -29182, -27024, -26004, -22271, -19733, -15463, 
    -10367, -6375, -2901, 1033, 6145, 11609, 13676, 18727, 22682, 23624, 
    26148, 27091, 30086, 31332, 31995, 31440, 28483, 28455, 24726, 22058, 
    20360, 16848, 10564, 8008, 4165, -265, -5492, -10755, -14056, -18659, 
    -21273, -23882, -27641, -28581, -30174, -30694, -31007, -30149, -29790, 
    -27432, -27263, -21452, -18659, -15577, -12137, -7632, -2318, -1, 5648, 
    9956, 14713, 17191, 21269, 25386, 25428, 27253, 29171, 31184, 30012, 
    30156, 29481, 28393, 25227, 21710, 19641, 15928, 11862, 8445, 4089, 
    -2066, -5049, -8093, -13059, -18021, -19317, -23021, -26700, -29530, 
    -31370, -30194, -31970, -30945, -29191, -28424, -25549, -22402, -19624, 
    -15730, -12458, -8701, -2823, -627, 5137, 8092, 12881, 16151, 20009, 
    22705, 25440, 28836, 29339, 32129, 29836, 30831, 29955, 28670, 25458, 
    23702, 20198, 17038, 12398, 9245, 4280, 823, -5891, -10158, -12590, 
    -16851, -19323, -22710, -24330, -27819, -30150, -30178, -30579, -31384, 
    -29533, -26430, -25859, -23412, -20586, -16481, -11739, -10330, -4060, 
    -120, 3153, 8473, 13103, 15744, 19022, 23513, 26891, 28080, 29569, 28936, 
    29378, 28795, 29399, 27736, 26318, 23981, 20298, 16307, 12599, 8983, 
    4402, -1355, -5178, -7396, -14300, -16379, -18518, -24693, -25737, 
    -28478, -29694, -30494, -29567, -30728, -29770, -29043, -25824, -23501, 
    -21196, -17065, -13001, -10486, -4965, -1903, 4613, 9646, 13247, 17669, 
    19683, 22699, 26824, 27974, 30321, 28708, 29658, 30843, 30486, 28217, 
    26452, 24480, 20633, 17068, 14523, 10162, 5319, 1101, -2832, -6393, 
    -12590, -15777, -19825, -22699, -25250, -27069, -28676, -30406, -31248, 
    -31312, -30213, -29807, -25820, -24163, -19068, -16883, -14008, -9505, 
    -5357, -972, 3856, 7409, 10744, 14900, 19832, 23203, 23772, 26555, 29243, 
    31637, 30754, 30421, 29396, 29825, 26465, 24337, 20986, 17411, 12935, 
    8932, 4292, 119, -4143, -6612, -12527, -15832, -20371, -23391, -25673, 
    -28448, -30684, -29604, -31126, -29591, -29781, -28172, -26009, -23824, 
    -22099, -19449, -15487, -9890, -6125, -928, 4185, 7156, 12638, 15964, 
    18220, 21632, 26350, 26087, 29979, 30725, 29206, 30900, 30973, 29558, 
    26801, 24215, 22257, 16705, 13121, 9647, 5272, 2134, -3409, -6741, 
    -11276, -15364, -17967, -21136, -25111, -27129, -28833, -29715, -31428, 
    -29062, -29563, -28579, -25745, -24441, -22402, -17363, -14203, -10776, 
    -5992, -2375, 1879, 6589, 12096, 14269, 18488, 22552, 24421, 28158, 
    29133, 30431, 30474, 31431, 30339, 29179, 27104, 24315, 22160, 17735, 
    15168, 9738, 5367, 1554, -3054, -7660, -11169, -15871, -18080, -21858, 
    -23673, -27009, -29729, -30464, -29854, -30354, -29105, -28355, -27400, 
    -23058, -21240, -18593, -16040, -10638, -6535, -1508, 2814, 7078, 11068, 
    13329, 19021, 21191, 23911, 26350, 28009, 29880, 29834, 29838, 28992, 
    28620, 27010, 23848, 22105, 16704, 15260, 11343, 6094, 2344, -189, -6177, 
    -9897, -15030, -17964, -20742, -24867, -26596, -27421, -30193, -30184, 
    -29571, -30941, -27468, -27061, -25198, -21430, -18837, -14530, -12449, 
    -7982, -2787, 1630, 7070, 9443, 14577, 17892, 22590, 24772, 27572, 30252, 
    30819, 29692, 30802, 31005, 28599, 26476, 23895, 23871, 19936, 16202, 
    11050, 8595, 4119, -867, -6727, -8707, -14259, -18495, -21223, -23863, 
    -26086, -30274, -28832, -30063, -30719, -32030, -31021, -27069, -23786, 
    -22165, -19048, -14585, -11813, -7437, -2944, 1249, 4708, 11185, 14390, 
    17309, 21387, 23736, 26260, 29296, 29562, 29220, 30290, 30948, 30825, 
    27552, 25916, 21910, 19308, 16071, 12482, 8368, 3333, 145, -6354, -9392, 
    -15136, -18973, -21428, -23443, -27192, -28091, -31345, -30629, -31432, 
    -29243, -28863, -27707, -25177, -22096, -20141, -15906, -12809, -7306, 
    -2700, 802, 5805, 8632, 12321, 17861, 20000, 24355, 24733, 28356, 29820, 
    30984, 30562, 30494, 27990, 27893, 25870, 22369, 19642, 15829, 13141, 
    8948, 3661, 266, -5446, -9861, -12383, -16350, -20532, -25189, -25632, 
    -27776, -28334, -31111, -30540, -31221, -28220, -27105, -25163, -22888, 
    -20122, -16307, -13206, -8658, -3409, -1378, 6061, 9039, 12985, 18110, 
    21041, 23216, 25879, 28848, 29778, 29613, 29438, 29244, 30203, 29345, 
    25334, 22759, 20942, 16721, 12137, 7900, 4546, 583, -5362, -9878, -12626, 
    -16542, -19794, -23081, -25524, -27233, -29620, -31655, -32247, -29847, 
    -30395, -27491, -26254, -23578, -19476, -15521, -11571, -8971, -4175, 
    573, 3897, 8182, 13866, 15629, 19263, 22909, 25307, 28030, 30065, 31055, 
    32402, 30659, 28744, 28543, 26617, 22241, 19551, 17199, 13526, 9509, 
    4792, -630, -4576, -7602, -12821, -17119, -20148, -22863, -25094, -26728, 
    -30267, -30825, -31355, -30555, -29360, -26360, -26324, -25094, -19275, 
    -17564, -12887, -8118, -5316, -1238, 3084, 10112, 12083, 17299, 20212, 
    23103, 24448, 27826, 29582, 30555, 29230, 31908, 31252, 28412, 25414, 
    23636, 22439, 17121, 13654, 7871, 5685, 673, -3103, -8235, -12194, 
    -15727, -20324, -23019, -24249, -29053, -29585, -31351, -32023, -30632, 
    -30274, -27588, -27133, -23636, -19760, -16068, -15239, -9030, -6450, 
    -1684, 3206, 7549, 12595, 16044, 19538, 22812, 25630, 27622, 28616, 
    29003, 30386, 30766, 28385, 27775, 26310, 23305, 20197, 17590, 13250, 
    10275, 5835, 1019, -3515, -7934, -11085, -15123, -19312, -21493, -24867, 
    -26560, -29225, -30829, -30067, -29095, -29602, -29677, -27839, -23951, 
    -19415, -18999, -12541, -11058, -5095, -984, 3291, 6495, 10670, 15697, 
    18734, 22168, 26696, 28214, 29520, 29364, 31026, 30049, 29987, 29967, 
    26702, 23853, 21729, 18360, 13487, 9599, 5269, 908, -2727, -7327, -12194, 
    -15069, -17386, -20962, -25749, -27588, -27886, -30386, -30748, -31229, 
    -30703, -28123, -26729, -25901, -20365, -17478, -13280, -9650, -5457, 
    -2204, 2940, 5664, 10785, 14558, 19028, 21779, 24848, 27516, 29128, 
    30687, 30863, 31865, 28833, 27567, 27444, 24975, 20436, 18623, 15458, 
    10605, 7077, 2220, -1761, -8038, -10677, -14450, -17609, -20987, -23867, 
    -28917, -28159, -30235, -30110, -30304, -30770, -27964, -27339, -23166, 
    -20633, -17290, -15053, -10129, -6326, -1471, 1101, 6514, 10063, 15664, 
    18653, 23519, 23887, 27447, 28203, 29391, 30253, 31376, 29982, 29473, 
    27453, 23533, 22116, 17359, 15269, 9142, 6935, 3187, -2387, -5809, -9979, 
    -13874, -18092, -20360, -23892, -25667, -28315, -31541, -29839, -30567, 
    -29609, -29620, -27581, -25774, -22459, -18395, -14576, -12793, -6952, 
    -3927, 2082, 7250, 10368, 13271, 17426, 21138, 25421, 26711, 28706, 
    29787, 29641, 31446, 31057, 29128, 27561, 24804, 21822, 18962, 14200, 
    11639, 7372, 2607, -2311, -5493, -10950, -14852, -18368, -21896, -22930, 
    -27477, -28177, -30992, -29306, -29921, -31147, -28812, -26809, -24784, 
    -21652, -18261, -14288, -10167, -7580, -3240, 1651, 6063, 10503, 13813, 
    18880, 21473, 23470, 26704, 28649, 30793, 30508, 29599, 31186, 28665, 
    28022, 26041, 23035, 19020, 14767, 11388, 8271, 3552, -571, -5415, 
    -11153, -13668, -16519, -20201, -22962, -26633, -29658, -31430, -31666, 
    -30290, -31817, -28632, -27590, -25504, -22699, -19557, -15837, -11954, 
    -8524, -4372, -114, 3873, 9541, 13634, 18329, 22419, 23869, 25271, 28130, 
    29656, 29962, 29755, 29739, 29502, 27507, 24805, 21313, 20634, 16307, 
    12899, 8507, 3003, -1462, -3626, -10507, -13197, -16511, -21042, -22383, 
    -26877, -28055, -29613, -31048, -30999, -30806, -28789, -28201, -24814, 
    -23252, -18905, -16000, -12157, -7778, -4066, -108, 6594, 9711, 13157, 
    15680, 21495, 22345, 25537, 29038, 29073, 30424, 30163, 30413, 30221, 
    27432, 24866, 22489, 19216, 15906, 11102, 9076, 4316, 478, -4627, -9624, 
    -13838, -16575, -20368, -23580, -26099, -29102, -27804, -29346, -30378, 
    -29132, -30865, -27305, -25915, -22450, -19433, -16671, -13056, -8838, 
    -4859, 244, 5525, 9063, 13059, 16128, 20069, 22941, 24797, 26503, 30216, 
    29376, 30278, 31238, 29822, 29967, 26094, 23420, 21738, 16608, 14724, 
    7928, 3937, 16, -5197, -8650, -12715, -17510, -18814, -23500, -24755, 
    -27639, -28363, -30202, -29833, -31141, -30465, -27141, -26349, -23871, 
    -20506, -17897, -12749, -9574, -4321, 515, 3925, 9191, 11935, 16752, 
    19289, 22902, 26258, 29021, 29168, 29997, 29374, 31550, 30457, 27782, 
    27427, 23364, 20827, 17655, 12852, 9899, 4838, -839, -4038, -6570, 
    -13070, -15938, -19200, -22209, -27008, -27578, -28784, -31516, -30606, 
    -30952, -29300, -27501, -25930, -23427, -19574, -17150, -14533, -9080, 
    -4200, -1433, 2241, 6932, 11219, 15926, 19433, 22360, 25028, 27558, 
    28426, 29953, 32457, 30761, 29975, 28300, 25510, 25148, 20828, 15899, 
    12914, 8922, 4209, 1269, -4131, -8795, -12779, -15512, -18672, -22194, 
    -24857, -27364, -30880, -30109, -31022, -30483, -30244, -27967, -27416, 
    -24965, -20376, -16939, -13491, -11114, -4531, -999, 2345, 6949, 11867, 
    16456, 20720, 21844, 26645, 28287, 28453, 31064, 30415, 30481, 29539, 
    28877, 28355, 24191, 22571, 18395, 14007, 10584, 5906, 820, -3910, -8007, 
    -10825, -15310, -18839, -22342, -25527, -27322, -29030, -30759, -32003, 
    -30740, -30935, -28679, -27911, -23304, -20224, -19256, -14611, -10541, 
    -5978, -2184, 1510, 6630, 10547, 14586, 19738, 21273, 26272, 26559, 
    30447, 30995, 32169, 30344, 29076, 28401, 27739, 24250, 21272, 19506, 
    14776, 11410, 5246, 1815, -2535, -6317, -10381, -14242, -18888, -22121, 
    -24893, -27754, -28087, -30451, -31414, -29448, -29547, -29656, -26329, 
    -24688, -23037, -18568, -14509, -11363, -6844, -2340, 1486, 7694, 10876, 
    15744, 18991, 22335, 24316, 27020, 28872, 30020, 30243, 31134, 31971, 
    30671, 27455, 23530, 21418, 18359, 14924, 10753, 6317, 2680, -1754, 
    -6805, -10721, -14028, -18914, -20399, -24185, -27524, -28716, -30328, 
    -30533, -30802, -29074, -28651, -27452, -24963, -21789, -18641, -14709, 
    -12177, -6403, -2661, 1541, 5954, 10885, 12883, 18479, 20669, 24069, 
    28260, 28792, 29515, 29999, 29618, 29843, 29750, 26380, 25557, 22030, 
    18310, 16279, 12414, 7717, 3991, -2431, -5553, -9342, -14850, -17898, 
    -22547, -23826, -27014, -26852, -30636, -31311, -32401, -30451, -29217, 
    -28964, -25178, -22231, -18723, -14028, -11575, -8703, -3608, 703, 3888, 
    11336, 12908, 18437, 22822, 24991, 26407, 27720, 29968, 29784, 30418, 
    31527, 29858, 26328, 26274, 22809, 20104, 15566, 12238, 7261, 4055, 
    -1551, -5533, -10358, -13469, -18002, -22741, -23607, -25758, -27205, 
    -30046, -30216, -30144, -30056, -27874, -26499, -26279, -24352, -19678, 
    -17017, -12074, -7435, -2769, -451, 5272, 9978, 12098, 17722, 19978, 
    23266, 26022, 28087, 28502, 31706, 32115, 31321, 27831, 27749, 25892, 
    22027, 18409, 16152, 10435, 8116, 3723, -1383, -3776, -8185, -13477, 
    -17696, -19800, -23333, -24410, -28139, -29328, -30070, -31406, -31293, 
    -28979, -26905, -26243, -23765, -20856, -15653, -12866, -8202, -4875, 
    1493, 3448, 8906, 13798, 17525, 21417, 23542, 25225, 27843, 29531, 30529, 
    30360, 31177, 28137, 28837, 26653, 23645, 21230, 17920, 11796, 8923, 
    4888, 326, -4302, -8570, -12691, -17023, -19911, -23966, -25294, -28387, 
    -29714, -30979, -31750, -29450, -28974, -27046, -25467, -23291, -19428, 
    -16231, -12786, -8522, -5063 ;
}
